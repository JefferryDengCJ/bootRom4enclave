/* Copyright 2018 ETH Zurich and University of Bologna.
 * Copyright and related rights are licensed under the Solderpad Hardware
 * License, Version 0.51 (the "License"); you may not use this file except in
 * compliance with the License.  You may obtain a copy of the License at
 * http://solderpad.org/licenses/SHL-0.51. Unless required by applicable law
 * or agreed to in writing, software, hardware and materials distributed under
 * this License is distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
 * CONDITIONS OF ANY KIND, either express or implied. See the License for the
 * specific language governing permissions and limitations under the License.
 *
 * File: $filename.v
 *
 * Description: Auto-generated bootrom
 */

// Auto-generated code
module bootrom_64 (
   input  logic         clk_i,
   input  logic         req_i,
   input  logic [63:0]  addr_i,
   output logic [63:0]  rdata_o
);
    localparam int RomSize = 7822;

    const logic [RomSize-1:0][63:0] mem = {
        64'h00003070_32635f30,
        64'h7032645f_30703266,
        64'h5f307032_615f3070,
        64'h326d5f30_70326934,
        64'h36767205_10040000,
        64'h002a0100_76637369,
        64'h72000000_34418082,
        64'hff87b503_0200c7b7,
        64'h8082e388_020047b7,
        64'h953eff87_b7830200,
        64'hc7b70030_7032635f,
        64'h30703264_5f307032,
        64'h665f3070_32615f30,
        64'h70326d5f_30703269,
        64'h34367672_05100400,
        64'h00002a01_00766373,
        64'h69720000_00344100,
        64'h46454443_42413938,
        64'h37363534_33323130,
        64'hb7bd4805_00f58023,
        64'h40d006bb_02d00793,
        64'hf606dee3_80826105,
        64'hfef816e3_00d700a3,
        64'hfec78fa3_177d0785,
        64'h0007c683_00074603,
        64'h9836972a_00b507b3,
        64'h9281982e_8f0d1682,
        64'h00150813_9f2d9e8d,
        64'h02b64a63_0017b593,
        64'hfd378793_4017569b,
        64'h40175613_00054783,
        64'h00080023_982afcc3,
        64'h7ee3fef8_8fa302c6,
        64'hd6bbfe87_c783978a,
        64'h02078793_93811782,
        64'h28058742_0006831b,
        64'h088502c6_f7bb0105,
        64'h08b32601_48012681,
        64'h08f60463_852e86aa,
        64'h47a9e83a_00f10c23,
        64'he4421101_0107c783,
        64'h67980007_b8030be7,
        64'h87930000_07978082,
        64'h8082fec7_ede3fee7,
        64'hae230791_87aafec5,
        64'h77e39f3d_0107179b,
        64'h9f2d0085_971b0ff5,
        64'hf5938082_fef61de3,
        64'hfeb78fa3_078502c5,
        64'h796387aa_0ff5f593,
        64'hcf81962a_8b8d00c5,
        64'h67b38082_fed59ae3,
        64'hfee78fa3_07850585,
        64'h0005c703_fec7fae3,
        64'h96ae40f6_06b3962a,
        64'h87aa8082_00c7ea63,
        64'h96ae40f6_06b395ba,
        64'h962a00e5_07b30711,
        64'h9b71ffc6_0713ff07,
        64'hebe3fed7_ae230711,
        64'h07914314_872e87aa,
        64'h03057963_982affd6,
        64'h0813ef8d_8b8d00b5,
        64'h67b3000b_0a010800,
        64'h30703263_5f307032,
        64'h645f3070_32665f30,
        64'h7032615f_3070326d,
        64'h5f307032_69343676,
        64'h72051004_0000002e,
        64'h01007663_73697200,
        64'h00003841_00000040,
        64'h00000020_001ff000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_000a2d2d,
        64'h2d2d2d2d_2d2d2d2d,
        64'h2d2d2d2d_2d2d2073,
        64'h00000000_0000006d,
        64'h00000000_3a207473,
        64'h6f632065_6d69742d,
        64'h2d2d2d2d_2d2d2d0a,
        64'h000a0d72_6f727245,
        64'h20647261_43204453,
        64'h00000000_00000000,
        64'h37323a33_313a3332,
        64'h00000000_002d2d2d,
        64'h00000000_00343230,
        64'h32203331_206e614a,
        64'h00000000_00203a74,
        64'h61206465_6c69706d,
        64'h6f632c20_6576616c,
        64'h636e6520_656e6f74,
        64'h7379656b_20726f46,
        64'h00000000_00000a0d,
        64'h30303176_2c646c72,
        64'h6f57206f_6c6c6548,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h4c0b2769_4aa850cb,
        64'h462bdcd7_17dd6425,
        64'hf31f7c6f_9688a5ba,
        64'h83851701_ffd4aa0f,
        64'h4a0eaa51_3472a806,
        64'hec89165a_833251ee,
        64'h60b92f85_29dcaec6,
        64'hd1d96021_b69a6a57,
        64'h73706c82_d7e713db,
        64'h04d8ba45_f6f5b454,
        64'hc91e7a5e_c9ab6306,
        64'h3aface8c_4799a040,
        64'h0000bf29_00a4d4bf,
        64'h10ef1ba5_05130000,
        64'h05178082_61797a1a,
        64'h79ba795a_74fa641e,
        64'h60be2d40_00ef4581,
        64'h4605854a_c1cff0ef,
        64'h06000613_0a040513,
        64'h85a686ce_874a2900,
        64'h00ef0128_02000613,
        64'h85d229c0_00ef8526,
        64'h04000613_85a2e28f,
        64'hd0ef8552_04040593,
        64'h86260804_0a13aaff,
        64'hf0ef8526_01aca59f,
        64'hf0ef01a8_85a24605,
        64'ha63ff0ef_01a84605,
        64'h85caa43f_f0ef01a8,
        64'h04000593_ad5ff0ef,
        64'h852201ac_10040413,
        64'ha83ff0ef_00000417,
        64'h01a805fe_45852b67,
        64'he6030000_0797a6ff,
        64'hf0ef01a8_04000593,
        64'he8afd0ef_854e85ca,
        64'h86260409_09930ce9,
        64'h09130000_0917fec7,
        64'h98e30685_278500e6,
        64'h8023fac7_071bfdd7,
        64'hc7130200_06134781,
        64'h86a6e2ff_10ef2ce5,
        64'h05130000_0517e3bf,
        64'h10ef0028_3f2000ef,
        64'h854a002c_4629fe84,
        64'h9de30421_00043023,
        64'he55f10ef_03397933,
        64'h2f050513_00000517,
        64'he65f10ef_002841c0,
        64'h00ef2501_002c4629,
        64'h03395533_03c00993,
        64'he7df10ef_2fc50513,
        64'h00000517_fef49de3,
        64'h07a10007_b02387a2,
        64'h00a40020_14041363,
        64'he39f20ef_34078aa3,
        64'h00000797_3647b903,
        64'h00000797_3667c503,
        64'h842a0000_079783bf,
        64'h20ef65a1_01f41513,
        64'he61f20ef_36078e23,
        64'h00000797_45013887,
        64'h83a30000_07973807,
        64'h89234405_00000797,
        64'he57f20ef_3a07b223,
        64'h00000797_30579073,
        64'hea678793_00000797,
        64'h3007a073_47a13047,
        64'ha0730800_07935c00,
        64'h00ef3cf7_3a236521,
        64'h00000717_87aa5e20,
        64'h00eff1ff_10efc265,
        64'h0513ffff_3517f2bf,
        64'h10ef38a5_05130000,
        64'h0517f37f_10ef38e5,
        64'h05130000_0517f43f,
        64'h10ef38a5_05130000,
        64'h0517f4ff_10ef36e5,
        64'h05130000_0517f5bf,
        64'h10ef3625_05130000,
        64'h0517f23f_10eff352,
        64'hf74efb4a_ff26e3a2,
        64'he7860805_05132005,
        64'h85937145_02faf537,
        64'h65f1f23f_206f4207,
        64'h8fa30000_07974467,
        64'hc5030000_0797f37f,
        64'h206f0141_44a78a23,
        64'h00000797_46e780a3,
        64'h60a24705_00000797,
        64'h64024607_88230ff4,
        64'h75130000_0797f35f,
        64'h20ef842a_e406e022,
        64'h1141b7e1_48878323,
        64'h00000797_f5bf20ef,
        64'hf79f206f_01414807,
        64'h8c230000_079760a2,
        64'h6402cb91_4a474503,
        64'h00000717_4ae7c783,
        64'h00000797_80820141,
        64'h640260a2_00f40663,
        64'h47854cf7_35230000,
        64'h07174ca7_3e230785,
        64'h00000717_4d574403,
        64'h00000717_4e47b783,
        64'h00000797_6f8000ef,
        64'h6ea000ef_e022e406,
        64'h65211141_fee79be3,
        64'h08000713_0ff7f793,
        64'h80820007_c3633420,
        64'h27f30000_30703263,
        64'h5f307032_645f3070,
        64'h32665f30_7032615f,
        64'h3070326d_5f307032,
        64'h69343676_72051004,
        64'h0000002a_01007663,
        64'h73697200_00003441,
        64'h00000001_00000006,
        64'h00000009_00000016,
        64'h0000000e_00000014,
        64'h00000002_0000000c,
        64'h0000000d_00000013,
        64'h00000017_0000000f,
        64'h00000004_00000018,
        64'h00000015_00000008,
        64'h00000010_00000005,
        64'h00000003_00000012,
        64'h00000011_0000000b,
        64'h00000007_0000000a,
        64'h0000002c_00000014,
        64'h0000003d_00000027,
        64'h00000012_0000003e,
        64'h0000002b_00000019,
        64'h00000008_00000038,
        64'h00000029_0000001b,
        64'h0000000e_00000002,
        64'h00000037_0000002d,
        64'h00000024_0000001c,
        64'h00000015_0000000f,
        64'h0000000a_00000006,
        64'h00000003_00000001,
        64'h80000000_80008008,
        64'h00000000_80000001,
        64'h80000000_00008080,
        64'h80000000_80008081,
        64'h80000000_8000000a,
        64'h00000000_0000800a,
        64'h80000000_00000080,
        64'h80000000_00008002,
        64'h80000000_00008003,
        64'h80000000_00008089,
        64'h80000000_0000008b,
        64'h00000000_8000808b,
        64'h00000000_8000000a,
        64'h00000000_80008009,
        64'h00000000_00000088,
        64'h00000000_0000008a,
        64'h80000000_00008009,
        64'h80000000_80008081,
        64'h00000000_80000001,
        64'h00000000_0000808b,
        64'h80000000_80008000,
        64'h80000000_0000808a,
        64'h00000000_00008082,
        64'h00000000_00000001,
        64'h00000000_0000bfd9,
        64'h4781bfe9_fb341ee3,
        64'h4781c83f_f0ef0028,
        64'h80826151_794e854a,
        64'h79ae74ee_641260b2,
        64'hf39ff0ef_c9be854a,
        64'h002cff34_11e30297,
        64'hd163f2e6_84238f2d,
        64'h04052785_00044583,
        64'hf286c703_002706b3,
        64'h0e078713_478100b4,
        64'h09b3c9a9_cba6cdb6,
        64'h0014949b_9c950640,
        64'h0493fee7_9de307a1,
        64'h0007b023_0998003c,
        64'h8932842a_f5cefda6,
        64'he606f9ca_e222716d,
        64'h80826105_450564a2,
        64'h644260e2_fed743e3,
        64'h0007871b_0d042683,
        64'h00d70023_078500f4,
        64'h87330007_468300f4,
        64'h07334781_02f05263,
        64'h0d042783_d2dff0ef,
        64'h842e00e7_8023f807,
        64'h4713852e_84aa0007,
        64'hc70300d7_002397ae,
        64'h37fd0066_c693ec06,
        64'he426e822_00074683,
        64'h972e1101_0cc5a783,
        64'h0c85a703_b7c5fc89,
        64'h13e34781_d6dff0ef,
        64'h85268082_61454505,
        64'h69a264e2_69420cf4,
        64'ha4237402_70a2fe89,
        64'h13e30137_de6300e6,
        64'h80238f2d_04052785,
        64'h0006c703_00044583,
        64'h00f486b3_00c58933,
        64'h842e0cc5_2983c60d,
        64'h84aa0c85_2783e44e,
        64'he84af022_f406ec26,
        64'h71798082_45050c05,
        64'h24230cf5_26230cb5,
        64'h28230017_979b9f8d,
        64'h06400793_fee79de3,
        64'h07a10007_b0230c85,
        64'h071387aa_80826179,
        64'h797a649e_643eedef,
        64'h9ce3e11c_8fb90f21,
        64'h000f3703_611cfbc4,
        64'h10e30283_03132415,
        64'hfcb710e3_fef2bc23,
        64'h00f3c7b3_8ff5e587,
        64'hb783978a_1b078793,
        64'h078efff6_c693e586,
        64'hb683968a_1b068693,
        64'h068e02c7_e7bb0004,
        64'h871b02a1_0002b383,
        64'h02c4e6bb_0027079b,
        64'h0017049b_4701829a,
        64'hff079be3_fed7bc23,
        64'h072107a1_6314871a,
        64'h003c4401_e43efc58,
        64'h9fe30391_e314631c,
        64'h8edd972a_0087d7b3,
        64'h00d796b3_070e40d0,
        64'h043b0291_0002a703,
        64'h0003a683_03010393,
        64'h09010293_651cfab4,
        64'h18e302a1_fef29ae3,
        64'hfce7bc23_8f350287,
        64'h87936398_8eb9e587,
        64'h3703970a_1b070713,
        64'h070e0076_e6b303f3,
        64'hd3930013_9693e586,
        64'hb383968a_1b068693,
        64'h068e02c7_673bf382,
        64'h87930003_841b0044,
        64'h071b02c3_e6bb0014,
        64'h039b4401_0c850293,
        64'hfeee90e3_06a10721,
        64'he29c0057_c7b30077,
        64'hc7b38fa1_8fa50a07,
        64'h32830787_33836b20,
        64'h7704631c_872a0034,
        64'h832a4e65_03010813,
        64'h88fa4595_46150285,
        64'h0e931b01_0f93f5be,
        64'hf1b6fd1a_ed16e91e,
        64'hedb2e9ae_e5c2e1c6,
        64'hf972f576_f17e0f01,
        64'h0f131787_37831707,
        64'h36831687_36031607,
        64'h3583f8ae_f0a2eca6,
        64'he8cae53e_e136fcb2,
        64'hf4fa1487_33031287,
        64'h32831207_33831587,
        64'h38031507_38831407,
        64'h3e031387_3e830e07,
        64'h3903e4ca_13073f83,
        64'h10073583_0d873903,
        64'he0ca7b60_77640d07,
        64'h3903fc4a_11873783,
        64'h11073683_0c873903,
        64'hf84a1087_36030f87,
        64'h3f030c07_3903fe67,
        64'h90e30206_86930207,
        64'h8793ee90_ea8c0106,
        64'hb4230116_b0236f90,
        64'h6b8c0087_b8030007,
        64'hb8830c07_03131994,
        64'h39478793_ff4ae3a6,
        64'he7a23947_87137145,
        64'h00000797_00003070,
        64'h32635f30_7032645f,
        64'h30703266_5f307032,
        64'h615f3070_326d5f30,
        64'h70326934_36767205,
        64'h10040000_002a0100,
        64'h76637369_72000000,
        64'h34418082_28010113,
        64'h45012581_39832601,
        64'h39032681_34832701,
        64'h34032781_30838082,
        64'h28010113_00153513,
        64'h25813983_26013903,
        64'h26813483_8d5d0107,
        64'h47b38d5d_0116c7b3,
        64'h27013403_8d5d2781,
        64'h30830066_47b38d5d,
        64'h01c5c7b3_8d5d01f4,
        64'h480301f1_47030105,
        64'h45338fd9_01e14683,
        64'h01e44883_8fd50117,
        64'h473301d1_460301d4,
        64'h43038fd1_0066c6b3,
        64'h01c14583_01c44e03,
        64'h8fcd01c6_463301b1,
        64'h450301b4_48038fc9,
        64'h0105c5b3_01a14703,
        64'h01a44883_8fd90115,
        64'h45330191_46830194,
        64'h43038fd5_00674733,
        64'h01814603_01844e03,
        64'h8fd101c6_c6b30171,
        64'h45830174_48038fcd,
        64'h01064633_01614503,
        64'h01644883_8fc90115,
        64'hc5b30151_47030154,
        64'h43038fd9_00654533,
        64'h01414683_01444e03,
        64'h8fd501c7_47330131,
        64'h46030134_48038fd1,
        64'h0106c6b3_01214583,
        64'h01244883_8fcd0116,
        64'h46330111_45030114,
        64'h43030104_4e038fc9,
        64'h01014703_0065c5b3,
        64'h8fd901c5_453300f1,
        64'h468300f4_48038fd5,
        64'h01074733_00e14603,
        64'h00e44883_8fd10116,
        64'hc6b300d1_458300d4,
        64'h43038fcd_00664633,
        64'h00c14503_00c44e03,
        64'h8fc901c5_c5b300b1,
        64'h470300b4_48038fd9,
        64'h01054533_00a14683,
        64'h00a44883_8fd50117,
        64'h47330091_46030094,
        64'h43038fd1_0066c6b3,
        64'h00814583_00844e03,
        64'h8fcd01c6_46330071,
        64'h45030074_48038fc9,
        64'h0105c5b3_00614703,
        64'h00644883_8fd90115,
        64'h45330054_43030051,
        64'h46830067_c7b38f35,
        64'h00414603_00444e03,
        64'h00314583_00344803,
        64'h00214503_00244883,
        64'h00114703_00014783,
        64'h00144683_00044303,
        64'hbe6f60ef_850a108c,
        64'he19f50ef_100c1088,
        64'h09b00204_06938f8f,
        64'he0ef1008_4ec000ef,
        64'h10081aac_496000ef,
        64'h1aa885ca_864e4a00,
        64'h00ef1aa8_02000613,
        64'h85a64ac0_00ef1aa8,
        64'h02000613_85a248e0,
        64'h00ef1aa8_04000593,
        64'h22051763_eb4f50ef,
        64'h84b689b2_26113c23,
        64'h25313c23_26913423,
        64'h85b609a8_892e842a,
        64'h27213023_26813823,
        64'hd8010113_80824501,
        64'h00e7f463_47fd03f5,
        64'h47030000_30703263,
        64'h5f307032_645f3070,
        64'h32665f30_7032615f,
        64'h3070326d_5f307032,
        64'h69343676_72051004,
        64'h0000002a_01007663,
        64'h73697200_00003441,
        64'h80822301_01132001,
        64'h3a032081_39832101,
        64'h39032181_34832201,
        64'h34032281_3083c33f,
        64'he0ef0204_0513002c,
        64'h862600b4_9cefe0ef,
        64'h00285c20_00ef0028,
        64'h122c56c0_00ef1228,
        64'h85ca864e_576000ef,
        64'h12280200_061385d2,
        64'h582000ef_12280200,
        64'h061385a2_564000ef,
        64'h12280400_0593c0ff,
        64'h50ef8522_012cc69f,
        64'h50ef0128_00aca18f,
        64'he0ef00a8_60c000ef,
        64'h00a8122c_5b6000ef,
        64'h122885ca_864e5c00,
        64'h00ef1228_02000613,
        64'h02048593_5a4000ef,
        64'h8a3689b2_21413023,
        64'h84ba2131_34232091,
        64'h3c232211_34230400,
        64'h05931228_892e842a,
        64'h21213823_22813023,
        64'hdd010113_00003070,
        64'h32635f30_7032645f,
        64'h30703266_5f307032,
        64'h615f3070_326d5f30,
        64'h70326934_36767205,
        64'h10040000_002a0100,
        64'h76637369_72000000,
        64'h34418082_613d6d9a,
        64'h6d3a6cda_6c7a7b9a,
        64'h7b3a7ada_7a7a699e,
        64'h693e64de_647e006c,
        64'h8fa3016c_8f23017c,
        64'h8ea301dc_8e2300bc,
        64'h8da301ec_8d2300fc,
        64'h8ca3018c_8c2301fc,
        64'h8ba300ec_8b2301cc,
        64'h8aa300ac_8a23005c,
        64'h892301ac_8823007c,
        64'h87a3010c_8723008c,
        64'h86a300dc_862301bc,
        64'h89a34113_53138599,
        64'h87ad8535_40785813,
        64'h40135b93_4037dc13,
        64'h01ebef33_01fc6fb3,
        64'h40555d93_40935b13,
        64'h01b46433_00259f13,
        64'h00579f93_410e5c13,
        64'h4137db93_00181d93,
        64'h770266e2_00ec88a3,
        64'h00dc85a3_8729011c,
        64'h83234027_5d1300cc,
        64'h822301a3_e3b3009c,
        64'h8523014c_8423012c,
        64'h83a3013c_82a366c2,
        64'h00dc84a3_40f85393,
        64'h00671d13_66a200db,
        64'h6eb3f076_408e5e93,
        64'h005ee2b3_00731693,
        64'h40e5db13_e4364127,
        64'h5e930035_129301d5,
        64'hf5b301de_7e3301d8,
        64'h7833931e_01d7f7b3,
        64'h4155d313_01d57533,
        64'h01d77733_95ea4157,
        64'hd593979a_415e5793,
        64'h9e5e4155_5e13e872,
        64'h955a4157_5513ec2a,
        64'h973e4158_5713983a,
        64'h972e8531_40455e13,
        64'h41455413_01c4e4b3,
        64'h00451e13_01d57533,
        64'h41555813_9542987a,
        64'h02870733_86a54016,
        64'hda134116_d49301c9,
        64'h69330076_9e1301d6,
        64'hf6b34156_d51396f2,
        64'h9e7e0387_0833015c,
        64'h81a3862d_4068d893,
        64'h40365a93_40e8d913,
        64'h0109e9b3_00289813,
        64'h01d8f8b3_4158d693,
        64'h03470e33_98c29816,
        64'h00ac8123_41365993,
        64'h646e00ae_65330056,
        64'h151301d6_76334156,
        64'h58939636_008506b3,
        64'h02d70833_010c80a3,
        64'h76a600dc_80234086,
        64'hd8134106_de1301d6,
        64'hf6b34156_d61302c7,
        64'h053396ee_01d3f3b3,
        64'h01d37333_664e0357,
        64'h06b34153_d71393ba,
        64'h01d67d33_41565393,
        64'h6726963a_41535613,
        64'h97468755_933640c3,
        64'h03330097_76330133,
        64'h07339342_986a01db,
        64'hfbb301db_7b3301d7,
        64'hf7b301d5_f5b3415b,
        64'hd6939bf2_415b5b93,
        64'h9e1e9d2a_03280833,
        64'h40c383b3_9b3a8e65,
        64'h41565313_4157db13,
        64'h97b64155_d693959a,
        64'h95b6038d_0d33961e,
        64'h750293aa_036585b3,
        64'h78e293c6_03250533,
        64'h415e5e13_038803b3,
        64'h40770733_009e73b3,
        64'h989effe0_04b70137,
        64'h0e339726_9772037d,
        64'h08b30010_09b79e4e,
        64'h03670733_01df7f33,
        64'h8a5e415f_53139f52,
        64'h00688f33_03850e33,
        64'h895a97ca_41e787b3,
        64'h01cf7f33_415f5493,
        64'h00c78f33_97fa0385,
        64'h88b39f26_036787b3,
        64'h99c60387_0f3301df,
        64'hffb36aae_415fda13,
        64'h9fd69ffa_037808b3,
        64'h99c60345_8fb301d2,
        64'hf2b34152_da9392d6,
        64'h41595913_6baa41f6,
        64'h86b301f9_7fb3ffe0,
        64'h0fb792fe_037d09b3,
        64'h94ce0375_82b39936,
        64'h6a2a0010_093796d2,
        64'h96ca0295_04b30366,
        64'h86b364aa_99a60378,
        64'h09b3994e_94960387,
        64'h89336b6e_934a4163,
        64'h033301cb_7b33415b,
        64'h5a1300c3_0b33036d,
        64'h02b39996_7ba69352,
        64'h037709b3_9a4e0386,
        64'h833301d4_74334154,
        64'h5a939456_941a0377,
        64'h8a3393d2_03658433,
        64'h92a24153_d3936a62,
        64'h414888b3_6baa01c3,
        64'hfa3300c8_83b398de,
        64'h98d20255_02b372a6,
        64'h4152da93_01d2fdb3,
        64'h036888b3_929e4159,
        64'h591378ca_411f0f33,
        64'h011978b3_ffe008b7,
        64'h997a0010_09379f46,
        64'h9f4a0355_82b39996,
        64'h03e68f33_033709b3,
        64'h6f2a947a_79a69a4e,
        64'h03680433_69c2994e,
        64'h035d8a33_9f220347,
        64'h89336aae_92d6032d,
        64'h0f337a26_036502b3,
        64'h405484b3_01c2f2b3,
        64'h4152db93_00c482b3,
        64'h94d29ffa_405f0f33,
        64'h01c2f2b3_4152d893,
        64'h00cf02b3_99960324,
        64'h84b39f46_036709b3,
        64'h03e68f33_74ca8926,
        64'h9aca7f26_98fa0358,
        64'h0ab384d6_92a60367,
        64'h88b3415f_df934113,
        64'h0333011f_f8b3ffe0,
        64'h08b79f46_035504b3,
        64'h9f9a0010_0fb7937e,
        64'h934e0357_0f330366,
        64'h8333999a_41e383b3,
        64'h01cf7f33_415f5f93,
        64'h00c38f33_01ef83b3,
        64'h035789b3_40740433,
        64'h01c3f3b3_9a4e4153,
        64'hda130346_8fb300c4,
        64'h03b379c2_00798433,
        64'h93a68ad2_93fe035b,
        64'h84b36b4e_036f8fb3,
        64'h93a66b86_6fa2997e,
        64'h6b6a408f_8fb301c4,
        64'h74334154_599300cf,
        64'h84339fa2_036b83b3,
        64'h41595913_407282b3,
        64'h01c973b3_00c28933,
        64'h92ce929e_035f8fb3,
        64'h6fa294fe_035903b3,
        64'h8bca6b0a_941e036b,
        64'h84b392a6_7b060369,
        64'h04339fa2_036b82b3,
        64'h69469396_7baa032b,
        64'h84336b6a_792294ca,
        64'h036383b3_73aa989e,
        64'h408888b3_01c47433,
        64'h41545993_036984b3,
        64'h00c88433_98a24153,
        64'hd3938bce_40930333,
        64'h01c3f4b3_00c303b3,
        64'h931e9326_035b8433,
        64'h7baa9fde_92a27bd2,
        64'h035b84b3_028b8433,
        64'h89de9926_03f98fb3,
        64'h7f8a0289_893398fe,
        64'h934a03fb_8fb36952,
        64'h92ca03f9_83336b0a,
        64'h74927406_7932989a,
        64'h6fea7bc6_63720269,
        64'h82b3405f_0f3301c2,
        64'hf2b34152_d39300cf,
        64'h02b37322_e49a9f1e,
        64'h406f8333_01237333,
        64'h41535593_937e0369,
        64'h88b3fc46_9fae4112,
        64'h88b30128_f8b34158,
        64'hdf939896_83460010,
        64'h08b792c6_03598f33,
        64'h63b2981e_41585813,
        64'h40650533_01c87333,
        64'h00c50833_957e951a,
        64'h028d02b3_ffe00937,
        64'h934a0285_0533975e,
        64'h875569ca_03898333,
        64'h650e8f89_01c77533,
        64'h00c78733_97fa97c2,
        64'h40eb8bb3_01c77733,
        64'h41575f93_00cb8733,
        64'h9b9a0287_07b3028b,
        64'h8bb3776a_40f705b3,
        64'h96ae01c7_f7b34157,
        64'hd69300c7_07b3973e,
        64'h977ef02a_40568533,
        64'h98aa01c2_f2b34152,
        64'hd89300c6_82b396c6,
        64'h96960284_8733983a,
        64'h02d486b3_74ca86a6,
        64'h9336038b_88334105,
        64'h85b301c8_78334158,
        64'h5f1300c5_883395fa,
        64'h03880333_9f9a028d,
        64'h85b392ae_038d8fb3,
        64'h977e025d_82b3680e,
        64'h96c27d8e_029d8733,
        64'h8d1901c7_77334157,
        64'h579300c5_07336d8e,
        64'h953e03b9_86b3ec3a,
        64'h8f1501c6_f6b34156,
        64'hd8939346_03850533,
        64'h00c706b3_973603b3,
        64'h0333754a_02570733,
        64'h9f2a84ee_774a9fba,
        64'h03848f33_95fa0259,
        64'h8fb3849a_029305b3,
        64'h97ae736a_969a03bf,
        64'h87b3953e_029f86b3,
        64'h9f3603bb_85337f8e,
        64'h98fe034b_8f3395aa,
        64'h025b88b3_937a0258,
        64'h85b397ae_03488333,
        64'h6daa951a_025d87b3,
        64'h78ea9fc6_029b8533,
        64'h95be029d_8fb372a6,
        64'h93160299_85b398fe,
        64'h034d8333_982e4158,
        64'h581375ae_8f0d01c8,
        64'h75b300c7_08339742,
        64'h034988b3_972e9746,
        64'h6a2e036a_05b39d1a,
        64'h64ce40a5_83b301c5,
        64'h75334155_531300c5,
        64'h853302a3_88b395a6,
        64'h971a0289_85b37506,
        64'h9f2ae82e_40b885b3,
        64'h01c5f5b3_4155df13,
        64'h03e70733_646e00c8,
        64'h85b398a2_98ae6d12,
        64'h6d8e7382_79ee7f22,
        64'h6762933a_035d05b3,
        64'h41585813_03330333,
        64'h97ae41e7_87b301c8,
        64'h7f3300c7_883397c2,
        64'h97fa03ba_08336342,
        64'h406f8fb3_01c37333,
        64'h41535593_00cf8333,
        64'h9f9a9fae_036387b3,
        64'h98c2035a_05b3972e,
        64'h6a6603ba_08b3798a,
        64'h9fc6033d_07337d62,
        64'h95ea03b3_8fb340d7,
        64'h86b301c6_f6b392ba,
        64'h4156d293_00c786b3,
        64'h979697b6_034585b3,
        64'h7382981e_035f86b3,
        64'h6fe2f87e_40df8fb3,
        64'h01c6f6b3_4156d413,
        64'h03640833_00cf86b3,
        64'h9fb6035a_06b39f36,
        64'h69a698c2_033f0f33,
        64'h6b0a6f62_41e70733,
        64'h01cf7f33_415f5313,
        64'h00c70f33_036f08b3,
        64'h97c6971a_03b787b3,
        64'h6f6293fa_03570733,
        64'h6b0a67c2_036783b3,
        64'h77029fba_67a29d3e,
        64'h03b40fb3_981e03a4,
        64'h0d3396fe_64060364,
        64'h083389da_033406b3,
        64'h933698c2_03b30333,
        64'h7b066442_8d0101c4,
        64'h74334154_52930368,
        64'h88b300c5_04336362,
        64'h951a78e2_9f460353,
        64'h03339722_63420333,
        64'h0f336346_406f0933,
        64'h012284b3_03648733,
        64'h97ba01c3_73334153,
        64'h529300cf_0333794e,
        64'h9f4a9f1a_02f487b3,
        64'h9f960333_033364a2,
        64'h636679a2_939a0334,
        64'h8fb377c2_96fe02f4,
        64'h83b3036f_8fb3981e,
        64'h6fc2957e_030a0833,
        64'h7a669752_03b48533,
        64'h77a27806_98c26dea,
        64'h74e202e4_8733942a,
        64'h033788b3_03b48433,
        64'h9f460347_8a3364c6,
        64'h92a6033f_0f33798a,
        64'h7f020334_02b3937a,
        64'h969669a6_03340333,
        64'h03b282b3_939a72e2,
        64'h798a9f96_033383b3,
        64'h6386981e_03640fb3,
        64'h79a27466_9522033f,
        64'h88337fc6_02a78533,
        64'h98fe6b0a_f5da7522,
        64'h40a80b33_01c57533,
        64'h41555913_00c80533,
        64'h984a0335_08b36562,
        64'h94aa03b8_893368e6,
        64'h01288f33_029584b3,
        64'h96fa0339_093384ca,
        64'h932669a6_033686b3,
        64'h76e679a2_92b60334,
        64'h84b393da_03b906b3,
        64'h7b72e25a_64a202d5,
        64'h83b39426_690666ca,
        64'hf94a4076_8b3301c3,
        64'hf3b3995a_4153d913,
        64'h00c683b3_7b4a0334,
        64'h043396da_969ef14e,
        64'h74467b0a_9fa20363,
        64'h83b303f5_8fb363e6,
        64'h981e7d86_6fc2957e,
        64'h03b80833_03a90533,
        64'h7da2886e_98c29f2a,
        64'h032588b3_93466922,
        64'h03390f33_92fa6906,
        64'h03690333_6b26006b,
        64'h04b30292_82b362a2,
        64'h7b2e9696_03630333,
        64'h634a03b5_86b3941a,
        64'h93b67d82_03ad8433,
        64'h9fa27de2_033d86b3,
        64'h74a29836_02990fb3,
        64'h6de2956e_03a906b3,
        64'h74c200d4_88b30365,
        64'h05339f46_02f586b3,
        64'hf1fe6946_fd4a6522,
        64'h40a68fb3_997e01c5,
        64'h75334155_5f93033f,
        64'h8f3300c6_8533796a,
        64'h96ca96aa_92fa03a5,
        64'h05336b26_f15a6fc6,
        64'h6566f9aa_41f50533,
        64'h01cfffb3_415fdb13,
        64'h03ab02b3_00c50fb3,
        64'h957e9316_6b62033b,
        64'h0fb3025f_82b36b66,
        64'h93da7fe6_798a947e,
        64'h033383b3_7f96987e,
        64'h02e40433_72c29d96,
        64'h03f40fb3_87a294be,
        64'h63c20275_82b36792,
        64'h969603a7_84b37fc2,
        64'h63c698fe_77c689be,
        64'h029982b3_e19e02f4,
        64'h0fb374c2_93a6742a,
        64'h9522405f_8bb301c2,
        64'hf2b34152_d49300cf,
        64'h82b39f96_72f69f96,
        64'h02fb8433_89de02e9,
        64'h82b39696_034b8fb3,
        64'h02e482b3_f97e7b82,
        64'h41f28fb3_034b86b3,
        64'h01cfffb3_415fd913,
        64'h00c28fb3_92a29f36,
        64'h76b66bc2_9f360375,
        64'h82b3034f_8f3389de,
        64'h951602e9_86b3987a,
        64'h6f76987a_02958533,
        64'h9daa79e2_9b4e6536,
        64'h00d50db3_034d8833,
        64'h02b989b3_67a66f56,
        64'h98fa64e2_651698aa,
        64'h029786b3_7fe6750e,
        64'hfdaa40d3_83b301c6,
        64'hf6b34156_d51300af,
        64'h833303ad_88b31efd,
        64'h00200eb7_7f4eea42,
        64'h00c386b3_02e90533,
        64'hf24674c2_6dca00dd,
        64'h843377c6_fa227dd6,
        64'h92ee8caa_034b83b3,
        64'hee666906_6be6008b,
        64'hf4330088_78330083,
        64'h78b3008e_fcb30058,
        64'h5813001b_db930073,
        64'h531303a3_86b3002e,
        64'hde93f636_019bebb3,
        64'h01e36333_01096833,
        64'h8ee18291_03620174,
        64'hebb303a2_82b37382,
        64'he61e6dd2_0bc201be,
        64'heeb304a2_018d9913,
        64'h79e20088_f3b30343,
        64'h8fb301d9_eeb301ff,
        64'h6f330f42_09a262c2,
        64'h7bca0058_68339b5e,
        64'h63a29b3e_0078e8b3,
        64'h011968b3_6bb2010b,
        64'h9893638e_00d3e6b3,
        64'h018c9393_0076e6b3,
        64'h01089693_87b60842,
        64'h09220172_e2b37b6e,
        64'h02a2010b_1e93016f,
        64'hefb3e2f6_0fa202f6,
        64'h86b30063_e3b303a2,
        64'h668600e6_c4839ea6,
        64'h0056cd83_0016c903,
        64'heeeefeca_00b6c383,
        64'h00c6c883_e69ee546,
        64'h0096cf03_0046c803,
        64'h0086cf83_0066c983,
        64'h77c20036_c28302e7,
        64'h8db300a6_c30300d6,
        64'hcc830026_cb830076,
        64'hcb035d18_0c130002,
        64'h1837008e_feb3fd42,
        64'h002ede93_03a303b3,
        64'h410f0833_01c87833,
        64'h41585913_00cf0833,
        64'h65380893_ffe00e37,
        64'hfff0c837_9f5a0010,
        64'h063702ec_84b377c6,
        64'h732af496_b6780293,
        64'hfe46e21a_f596faee,
        64'heda6eaca_f1f2000a,
        64'h08370038_d893e9c2,
        64'h02f98f33_01fb8db3,
        64'he5faea6e_d1880813,
        64'hc13f0f13_0078e8b3,
        64'h000a3f37_008f72b3,
        64'h00073837_0058e8b3,
        64'h934208a2_006f5f13,
        64'h02c269e6_00887833,
        64'h9dce0058_5813018f,
        64'h6f330183_9f1302ff,
        64'h8fb30136_c8830116,
        64'h0bb3e65e_0146c283,
        64'h0126c383_0083fab3,
        64'h664e9db2_68ee02fc,
        64'h83330833_04930074,
        64'hd913fdca_7dea662e,
        64'h6fe2fff5_933701f8,
        64'h6833006c_6c3301e3,
        64'h63330c42_08627f4a,
        64'h997a0322_77c26f2a,
        64'h01e4e4b3_01889493,
        64'h029609b3_6ccaf9be,
        64'h008cfe33_01ccecb3,
        64'h0116cc03_0199ecb3,
        64'h005f6f33_76620106,
        64'h6eb303ae_8bb30f42,
        64'h09a201b2_e2b302a2,
        64'h74c2010b_9c93009f,
        64'hefb30fc2_0174e4b3,
        64'h02f587b3_7ee601d3,
        64'he3b377c6_9b3e008d,
        64'h7d3304a2_7ea6f976,
        64'h0106c303_01e6cf03,
        64'h0196cf83_0176cb83,
        64'hf2e202eb_8b330166,
        64'hc98301d6_c2830186,
        64'hc4830156_ce0301f6,
        64'hc88301a6_c803e172,
        64'hf0c6f442_034c8c33,
        64'he196f126_008e7e33,
        64'h0088f8b3_8ce10006,
        64'hc2838796_00cc6633,
        64'h010d9c13_02ec0933,
        64'h002e5e13_0078d893,
        64'h00f6ce83_8085ed76,
        64'h0138e8b3_008efeb3,
        64'h005ede93_01d36eb3,
        64'h034f82b3_6c22018c,
        64'h1313f69a_08e201e9,
        64'he9b309c2_7b820622,
        64'h012eeeb3_7cc6007c,
        64'he3b303c2_026a8333,
        64'h0ca2018e_6e337342,
        64'h00837833_e5420079,
        64'h693301b6_c60301c6,
        64'hcd830922_6fe20016,
        64'h4c830056_4c036ac2,
        64'h00435313_034a8833,
        64'h01081e93_01d36333,
        64'h03620064_e4b3017e,
        64'heeb30ec2_011bebb3,
        64'h6ac6e496_01caee33,
        64'h00364903_00964983,
        64'h00464803_00264383,
        64'h00385593_0e420aa2,
        64'h00b86833_01cf6f33,
        64'hf53ef8ee_e5caecce,
        64'he462008f_f2b30f22,
        64'h008cfdb3_006fdf93,
        64'h008d9b93_0082f7b3,
        64'h0079d993_edbe0022,
        64'hd29302e9_0933005c,
        64'hdc93019b_ecb30066,
        64'h4a830076_4e03e956,
        64'he8f2008a_fab3008e,
        64'h7e33007e_5e1302eb,
        64'h07b300f2_e2b38f61,
        64'h7966012d_6d336b42,
        64'he9da8309_77a27906,
        64'h01096833_09220842,
        64'hfd3e690e_682e0343,
        64'h8b33009b_64b304c2,
        64'h0b2273e2_01f3efb3,
        64'h01859393_007fefb3,
        64'h64a66b4a_0054e2b3,
        64'h016aeab3_01091f93,
        64'h008f9493_65ea7b46,
        64'h034587b3_01ab6d33,
        64'hf83e796a_0d420129,
        64'he9b30b22_8fe1007a,
        64'h5a138395_09e26586,
        64'h0085fc33_0183e3b3,
        64'h03a28191_6c26010c,
        64'h12930182_9b93017c,
        64'hecb30cc2_6c2272a2,
        64'h015c6ab3_005a6a33,
        64'hf04200a6_488300c6,
        64'h4e83ec46_e8760086,
        64'h4f0300d6_4303fc7a,
        64'hfc9a6b4e_e0a60169,
        64'h69337d42_73ca79aa,
        64'h6f8a00b6_4d830942,
        64'h003f5f13_7ce6008f,
        64'hf333010c_9a930083,
        64'h74b3008a_9c138fc5,
        64'h01876733_00887833,
        64'h0088f8b3_008efeb3,
        64'h019bebb3_00285813,
        64'h0058d893_0ba2013e,
        64'heeb3007f_6f33006f,
        64'hdf93018c_14930013,
        64'h53138fc5_147d0020,
        64'h043707c2_01841a13,
        64'h01a86833_01bf6f33,
        64'h01436333_6a860f22,
        64'h015eeeb3_790a0dc2,
        64'h012b6b33_6cc60b22,
        64'h0ea279e2_63c200b9,
        64'he5b3007e_6e336be6,
        64'h0ac2f0de_6d620e62,
        64'h011d68b3_018a1993,
        64'h646e0135_e5b30082,
        64'he2b37902_02c2012f,
        64'hefb30d62_01946433,
        64'h01c9e9b3_04220156,
        64'h4b8309a2_e95e6a2a,
        64'h0143e3b3_03c200e6,
        64'h4b83ed5e_6f4a6d62,
        64'h018f1f93_01a8e8b3,
        64'h01f36333_01e64283,
        64'h01964783_01d64403,
        64'h01a64c03_08c20322,
        64'h015d6d33_0d220126,
        64'h4b8300eb_e733010c,
        64'h97138cd9_6f4201e9,
        64'h69337742_00e86833,
        64'h09420ba2_676a0107,
        64'h159300ba_6a3304a2,
        64'h770665a2_e1bae5ae,
        64'h08220136_47030146,
        64'h4583e4ba_fd2e0a22,
        64'h00f64703_01164583,
        64'hed3a0105_97130107,
        64'h1f9300ef_6f33e9fe,
        64'h7582f92e_01664f83,
        64'hf87e0106_4583edae,
        64'h0f220176_4f8301f6,
        64'h458301b6_4b830186,
        64'h4483f4a6_f52ef122,
        64'hfc16e962_fcfe01c6,
        64'h4c8301f5_c5830115,
        64'hc9030095_c383f0ca,
        64'he11e0165_ce8300e5,
        64'hc303ecf6_e09a01d5,
        64'hcb0301b5_c8030195,
        64'hc8830145_cd8300b5,
        64'hc9830085_ca030006,
        64'h448301e5_c4030155,
        64'hc2830135_cc030045,
        64'hcf8300c5_c9030065,
        64'hc3830035_ce830015,
        64'hc303f8c6_0185cd03,
        64'h0105cf03_0175ca83,
        64'h00a5ce03_00f5c703,
        64'hf042ec26_e822e552,
        64'he43af43e_e8e60005,
        64'hc88301c5_c80301a5,
        64'hc4830125_c40300d5,
        64'hca030075_c7030055,
        64'hc7830025_cc83e76a,
        64'heb66fb56_ff52eba6,
        64'hefa2e36e_ef62f35e,
        64'hf75ae3ce_e7ca7105,
        64'h80826119_7d927d32,
        64'h7cd27c72_6b966b36,
        64'h6ad66a76_79967936,
        64'h74d601c5_0fa301e5,
        64'h0e2300b5_0da301f5,
        64'h0d2300f5_0ca30055,
        64'h0ba301d5_0aa30105,
        64'h0a230075_092300e5,
        64'h08a30165_0f230175,
        64'h0ea30185_0c230195,
        64'h0b2301b5_09a301a5,
        64'h0823411e_5e138599,
        64'h87ad40d8_58138729,
        64'h409e5b13_401e5b93,
        64'h01eb6f33_01fbefb3,
        64'h4037dc13_408edc93,
        64'h005c62b3_007ce3b3,
        64'h40585d93_40275d13,
        64'h74760085_07a3007e,
        64'h1f130025_9f930057,
        64'h9293410e_dc130038,
        64'h139340e5_db134137,
        64'hdb934127_5c930115,
        64'h072300d5_06230065,
        64'h032300c5_02234078,
        64'hd8930095_06a30145,
        64'h04230125_03a30135,
        64'h02a30155_01a301a4,
        64'h643301e5_f5b301ee,
        64'hfeb301e8_783301e7,
        64'hf7b340f8_d41301b4,
        64'he4b30067_1d139e22,
        64'h4155de13_00189d93,
        64'h01e77733_66c200d5,
        64'h05a395e2_01e8f8b3,
        64'h4157d593_979666a2,
        64'h00d50523_415ed793,
        64'h9e9e4158_5e936682,
        64'h00d504a3_985e4157,
        64'h5813e442_e02e975a,
        64'h4158d713_e83a98be,
        64'h97fe8731_40475813,
        64'h41475493_0105e5b3,
        64'h00471813_01e77733,
        64'h41575893_974698a6,
        64'h03b787b3_86a54016,
        64'hda134116_d5930109,
        64'h69330076_981301e6,
        64'hf6b34156_d71396f2,
        64'h9e520317_88b34063,
        64'h5313862d_00b9e9b3,
        64'h40e35913_00231593,
        64'h01e37333_41535693,
        64'h933696ca_03c78e33,
        64'h40365a93_41365993,
        64'h00e50123_8f4d0056,
        64'h171301e6_76334156,
        64'h5313963a_96420267,
        64'h86b36822_010500a3,
        64'h00d50023_4086d813,
        64'h4106d593_01e6f6b3,
        64'h4156d713_02c78633,
        64'h96d601e4_743301ec,
        64'h7c3302d7_86b34154,
        64'h5793943e_01e2f2b3,
        64'h415c5413_77c29c3e,
        64'h4152dc13_97ba87d5,
        64'h92f64088_02b38c7d,
        64'h97c29816_92ae01e3,
        64'hf3b36a82_674295ba,
        64'h03b282b3_4153de93,
        64'h67620137_03b399d6,
        64'h41da8ab3_008efeb3,
        64'h415ed813_00fa8eb3,
        64'h9af6031c_85b39a9e,
        64'h03be8eb3_01ebfbb3,
        64'h93ea0312_8ab301eb,
        64'h7b3301ef_ffb3415b,
        64'hd7139bae_415b5b93,
        64'h9b3a415f_db139fe2,
        64'h9fc203cc_83b301e4,
        64'hf4b34154_dc1394e2,
        64'h017384b3_03bf8fb3,
        64'h4159d993_415585b3,
        64'h0089fab3_00f589b3,
        64'h95ce95d6_031f83b3,
        64'h9ada03b5_85b39b1e,
        64'h031e8ab3_97568f05,
        64'h8ce14154_d99300f7,
        64'h04b39726_03c283b3,
        64'h94ce03b7_07339b1e,
        64'h031584b3_01ea7a33,
        64'h415a5c13_9a629a26,
        64'h026c8b33_99da03cf,
        64'h8a337c82_9b6603ce,
        64'h89b3415a_da934148,
        64'h0833008a_fa3300f8,
        64'h0ab39856_02628b33,
        64'h98529a5a_03b80833,
        64'h01e97933_41595c13,
        64'h99620317_0a337de2,
        64'h01b98933_026f89b3,
        64'h01390cb3_9bd2419b,
        64'h8bb3008c_fcb3415c,
        64'hda939b56_02c90933,
        64'h00fb8cb3_9be603c5,
        64'h8b339cda_03180bb3,
        64'h7902415b_dc13e44a,
        64'h01ebf933_9be29bca,
        64'h03c70cb3_02cf8bb3,
        64'h9ade9d66_415cdc93,
        64'h7d2241a3_83b3008c,
        64'hfd3300f3_8cb393ea,
        64'h93e6026e_8ab3e056,
        64'h01eafab3_415adc13,
        64'h9ae202c3_83b3415a,
        64'h5a136382_407484b3,
        64'h008a73b3_00f48a33,
        64'h94d2949e_02df8c33,
        64'h9b6203c8_04b39ba6,
        64'h02658b33_9cda02c2,
        64'h8bb37b26_93da02db,
        64'h8cb30267_03b3949e,
        64'h6ba29c5e_02dc84b3,
        64'h63a64079_89b30083,
        64'hf3b34153_dd1300f9,
        64'h83b399ea_02ce8c33,
        64'h7c829be6_02d989b3,
        64'h00748db3_418383b3,
        64'h008c7c33_415c5a13,
        64'h00f38c33_93d202d2,
        64'h8bb36982_9b4e0268,
        64'h03b39a1e_02c58b33,
        64'h93ee02c7_0a3399da,
        64'h02d583b3_84d54149,
        64'h09330084_fa3300f9,
        64'h04b39952_992602de,
        64'h89b3407a_8ab30083,
        64'hf3b34153_da1300fa,
        64'h83b39a9e_02c80933,
        64'h94ca02d8_0ab3f862,
        64'he85263c6_40798c33,
        64'h0083f3b3_4153df93,
        64'h00f983b3_999e6906,
        64'h02d704b3_40990a33,
        64'h8ce14154_d99300f9,
        64'h04b3997e_6de692d2,
        64'h4152d293_409e8eb3,
        64'h0082f4b3_00fe82b3,
        64'h9ece9e96_03b48933,
        64'h7a4692ca_03ba8eb3,
        64'h7482794e_95f68f05,
        64'h85d50085_f4b300f7,
        64'h05b39726_974a031a,
        64'h02b34055_8eb30082,
        64'hf2b34152_d99300f5,
        64'h82b395ce_03b70733,
        64'h7b069876_674240e3,
        64'h83b38f61_41575813,
        64'h00f38733_93e203bb,
        64'h05b30058_03b3ec2e,
        64'h407705b3_9fae0083,
        64'hf3b34153_df9300f7,
        64'h03b3975e_971e03bf,
        64'h88337a42_414585b3,
        64'h008a7a33_415a5c13,
        64'h00f58a33_95e203cf,
        64'h87339942_031585b3,
        64'h6f8299fe_031b0833,
        64'h40ee8eb3_8f614157,
        64'h549300fe_87339eba,
        64'h031989b3_92c28ace,
        64'h03ba8eb3_01d483b3,
        64'h991e031a_82b303c9,
        64'h89337de2_9fee026a,
        64'h84b36582_6b62f416,
        64'hf4a601e9_7d337da6,
        64'h808d0069_591301b4,
        64'he4b303ca_0fb30164,
        64'he4b3012f_e9336aa2,
        64'h79a24152_82b3e4ce,
        64'h04a2018d_9f930b42,
        64'h01f96933_008afab3,
        64'h01e9f9b3_415adb93,
        64'h0019d993_00f28ab3,
        64'h92de7a42_00b9e9b3,
        64'h01ea7cb3_004a5a13,
        64'h013ce9b3_7dae014d,
        64'h6a3365a6_f0ae01ea,
        64'hf5b30262_82b3972e,
        64'h007ada93_62820135,
        64'h4483ecee_01e2fdb3,
        64'h010d9913_01091993,
        64'h013aeab3_012fefb3,
        64'h0fa20022_d293694e,
        64'h7d8e0189_1d13008d,
        64'h9c93031d_07339866,
        64'he0ba01e7_77336fee,
        64'h83156926_012a6a33,
        64'h010f9a13_6dae0149,
        64'he9b36f8e_018f9a93,
        64'h01f96933_008d9913,
        64'h01276733_7fca01f2,
        64'he2b303cd_0cb37dea,
        64'h010d9993_0092e2b3,
        64'h01099493_01849713,
        64'h9c3a0145_4b03985a,
        64'h5d188893_000218b7,
        64'h013a6a33_6f8601fa,
        64'h8eb303cc_0c33e8f6,
        64'h01ecfeb3_7daa93f6,
        64'h01bcecb3_01eefeb3,
        64'h69ea6486_001ede93,
        64'h02cd0ab3_009cecb3,
        64'h0ca26de6_008d9a13,
        64'h7c86f4e6_7d8a008d,
        64'h92930059_6933026a,
        64'h03b30103_99136dca,
        64'h6d4295ea_63aa0072,
        64'he2b30103_94937a42,
        64'h00849293_f9960032,
        64'hd29373e6_0152e2b3,
        64'h9b9e03cd_0d33648a,
        64'h0142e2b3_f8a64129,
        64'h84b302a2_01e4fcb3,
        64'h0a429fe6_8099026d,
        64'h0b3301ef_ffb30089,
        64'h7933ffe0_0437005f,
        64'hdf939822_7cc695e6,
        64'h653e0e13_fff0ce37,
        64'h02cc0bb3_975e976e,
        64'h6c226452_8cc10285,
        64'h42836d62_971601af,
        64'hefb30295_4a0393e2,
        64'h6df295ee_018a9493,
        64'h01e3f3b3_6d92986e,
        64'h01e77733_62b27dee,
        64'h01beeeb3_005a6eb3,
        64'h010b1293_02628bb3,
        64'h8c450442_830901e5,
        64'hf5b30164_e4b304a2,
        64'h02754a83_75a6f8ae,
        64'h02dc0c33_01e87833,
        64'h02654403_00785813,
        64'h02554483_0a226dc6,
        64'h01b3e3b3_0173e3b3,
        64'h62c202de_85b30182,
        64'h9f930235_4a0301fd,
        64'h6d330245_4b030d42,
        64'h6c42008c_13937d46,
        64'h010d1b93_026b8cb3,
        64'h01976733_01afefb3,
        64'h8f41b673_03136ee2,
        64'hf0767282_9eae4159,
        64'h5593f4ae_819100b2,
        64'he5b3000a_033700f9,
        64'h893372ce_f9ca018a,
        64'h99137c82_7c266ac6,
        64'h00bae5b3_010c1a93,
        64'hea56008c_9f93ec5a,
        64'h01eefeb3_005ede93,
        64'h007eeeb3_99fe0010,
        64'h07b70ee2_00f3e3b3,
        64'h02cb8ab3_ee5601ef,
        64'hffb303c2_014fefb3,
        64'h8fc50058_68330189,
        64'h18130102_e2b30125,
        64'he5b37ba2_02cb0ab3,
        64'h010b9293_01029413,
        64'h008a9593_00859713,
        64'h00efefb3_01049713,
        64'he23af822_02a54a03,
        64'h033a09b3_07a20058,
        64'h68330822_0fa202e5,
        64'h438302d5_4783e446,
        64'hfdf2e61e_02c40733,
        64'he83efc4e_08398993,
        64'h01e8f8b3_01e7f7b3,
        64'h0078d893_8391fff5,
        64'h99b78452_02d403b3,
        64'h02b54f83_02c54483,
        64'h01effb33_0068e8b3,
        64'h08e2e03a_01e77733,
        64'hf4220073_633302da,
        64'h0e33d186_06130007,
        64'h36378309_00165f93,
        64'h034201f7_e7b301e4,
        64'h7433c136_8693000a,
        64'h36b70066_d41301d7,
        64'h67330184_17938e41,
        64'h00ffefb3_1f7d0020,
        64'h0f370fc2_01c76733,
        64'h01e66633_0117e7b3,
        64'h07220622_07a20e42,
        64'h0f420335_430301c3,
        64'he3b303a2_02f54e83,
        64'h03754403_01d6e6b3,
        64'he8a206e2_03654f83,
        64'h009eeeb3_03454883,
        64'h0ec20305_47030385,
        64'h46030355_478301e4,
        64'he4b30315_4e030037,
        64'h5a1304a2_03254383,
        64'h01376733_02254403,
        64'h07620069_e9b309c2,
        64'h03b54e83_00d36333,
        64'h03954f03_032203a5,
        64'h448303f5_470303e5,
        64'h498303c5_468303d5,
        64'h43030215_4c03f1e2,
        64'h01d54803_f8ba01e5,
        64'h4b83f4be_edde0205,
        64'h4a83e5da_e1d6fd52,
        64'hf57af176_e972e51a,
        64'he146f0c2_01b54583,
        64'h01854c83_01654783,
        64'h01154c03_8dbe0195,
        64'h47030105_4b8300e5,
        64'h4b0300c5_4a8300b5,
        64'h4a030095_4f030085,
        64'h4e830065_4e030045,
        64'h43030035_48830015,
        64'h48030155_4783eca2,
        64'h01f54903_01c54283,
        64'h01754d03_f02ef5b2,
        64'he9b6e4ba_f97eed4e,
        64'he0befc9e_f26ef66a,
        64'hfa66fe62_e2dee6da,
        64'head6eed2_f6cafaa6,
        64'h00054403_fea201a5,
        64'h45830125_460300f5,
        64'h468300d5_470300a5,
        64'h4f830075_49830055,
        64'h47830025_4383f2ce,
        64'h71090000_30703263,
        64'h5f307032_645f3070,
        64'h32665f30_7032615f,
        64'h3070326d_5f307032,
        64'h69343676_72051004,
        64'h0000002a_01007663,
        64'h73697200_00003441,
        64'h80826129_74aa744a,
        64'h70eaa4bf_70ef8526,
        64'h858aaa5f_70ef850a,
        64'h00f40fa3_00e40023,
        64'h0407e793_9b6103f7,
        64'hf79385a2_00044703,
        64'h01f44783_4c8020ef,
        64'hfd06853e_02000593,
        64'h04000693_84aa862e,
        64'h842ef526_f92287b2,
        64'h71310000_30703263,
        64'h5f307032_645f3070,
        64'h32665f30_7032615f,
        64'h3070326d_5f307032,
        64'h69343676_72051004,
        64'h0000002a_01007663,
        64'h73697200_00003441,
        64'h003fbe44_01191df9,
        64'hff2be4a0_01d0e833,
        64'hffa497ba_ffae1238,
        64'h007bf8cb_fe8fdc75,
        64'h00e43411_fec84266,
        64'h0046d77c_018a44cc,
        64'h00a87df4_014646fe,
        64'h00c84e2a_ffffbb60,
        64'h008d9738_ff5a0358,
        64'hff24abd2_01c5342e,
        64'h0065cd7f_017f6bc2,
        64'h0014dc50_ffe3b7e7,
        64'hffedaa49_fe3170e6,
        64'hffbcb56d_006b17ef,
        64'h00eee291_fea975fc,
        64'h009c8891_0112c7df,
        64'hff3c9bc4_fe298e30,
        64'h00e1c52b_01c34e0c,
        64'h000519a0_01e3a4bb,
        64'hff120c9f_ff95d543,
        64'h002df576_00a6c315,
        64'hff0b1929_fe24e98d,
        64'hff5f0367_feb810bd,
        64'hff9d22ac_003ce8c2,
        64'h00c1eccc_feed3e33,
        64'hff13b297_fe2a74be,
        64'hff3c2ee8_ff7dbbd5,
        64'h003ad61f_01e3c28e,
        64'hff877821_ff55254d,
        64'h00abea98_fe10b0cc,
        64'hffc3c0a8_fecf0c81,
        64'h0063e4e4_01f9b77c,
        64'h00cbb03b_ff48af06,
        64'hff31734a_01dffd61,
        64'h00976319_fffd2add,
        64'hffc27e91_ffedcb29,
        64'h003527f1_01e044bf,
        64'hff909459_fe3e5800,
        64'h00452540_ff996c25,
        64'h006ff841_00aa63aa,
        64'h00b2cb17_01f54516,
        64'hff456cbf_fe4971bf,
        64'hff3473f5_fe26bccc,
        64'h002e208b_feec1105,
        64'h00b2faff_01022790,
        64'hff655d83_015b508f,
        64'h00b2e70c_006cf8dc,
        64'hffe73e23_00c239b9,
        64'hff25bd68_00818717,
        64'hff3243bd_ffd7c223,
        64'h00b35af4_fe3fb1db,
        64'h00ec7532_01212ff1,
        64'hff3a476b_ff5b3be1,
        64'hffa3f7ff_00614e3c,
        64'hff0ef83e_00e6bba0,
        64'hffa2b3bb_fed9bd41,
        64'h0023f077_fed38b79,
        64'h00dab979_01266898,
        64'h0071a7e8_fe02c065,
        64'hfff5913d_ff233f31,
        64'hff28e588_fe2c918a,
        64'h002a83d5_01a138ec,
        64'h003245da_fee7b78f,
        64'h0016c18b_ff090232,
        64'hff462410_01e32da9,
        64'h0006ac4b_015807e3,
        64'h0042e145_ff67b17d,
        64'hff2800ba_0075a74e,
        64'hff352aaa_ff8f94ee,
        64'h00e0de2d_ffeb54d5,
        64'h0048fa9b_fe3354bd,
        64'h00a1d107_00478eb0,
        64'h0061e23b_001d1286,
        64'h00d8183c_ff037389,
        64'h002479fe_fed266fd,
        64'hff567541_00f7f6b8,
        64'hff7c92e4_feb48a58,
        64'hff8460d4_0132d528,
        64'h00c504cc_ff5abc5a,
        64'h006f19a4_00fe3914,
        64'h00955d45_0042a9fb,
        64'h006a2a31_ff6c581a,
        64'h00691fab_00823871,
        64'h0096b210_01f2a145,
        64'h0026f5c8_fe04f676,
        64'hffaeea0a_00f89699,
        64'hff337997_0117ef27,
        64'hff1be527_ff0d28c9,
        64'hff397e6c_00fc722c,
        64'hffdffd5e_fef121ba,
        64'h00978600_fe4d50ac,
        64'h00276326_00ce3b79,
        64'h009ab0ab_00b81e05,
        64'h0022c43f_0102c998,
        64'hff4d3a50_fe8a35af,
        64'h00e4b8eb_00aa8c87,
        64'hffc84ea0_feb63eb6,
        64'h002b5e02_fe07dba2,
        64'h00d3dd32_fee8356b,
        64'hff25123f_fec8f53e,
        64'hffb14d74_013ff776,
        64'h003ab907_00e355cd,
        64'hffdcdef2_fea074fc,
        64'hff7046d5_01efe9e8,
        64'hff95c110_fe7b01a7,
        64'h007ee886_00aef40b,
        64'hff685f09_00cfc88d,
        64'hff54fa8e_00822707,
        64'hff79d225_01921400,
        64'h00ffaf6e_01be82f0,
        64'h003e8d85_00f3b1ca,
        64'h00d7eba5_fea7f9cc,
        64'hff808679_fef232fb,
        64'h0072267e_fe741a59,
        64'hff812d89_fe943dff,
        64'hff001506_01b1d2bc,
        64'h00280df7_ff9f2a62,
        64'h00dfb635_ffe72681,
        64'hffae0ed6_00b6cd21,
        64'h000ac3a3_00936a63,
        64'h00703e80_01a36371,
        64'h0086dfd7_0161694b,
        64'hff3afa05_0172b9a9,
        64'hfffabe5e_01ec3f97,
        64'hff196276_fe3b5f39,
        64'h003d8be7_00332ba5,
        64'h008a8851_0089a66a,
        64'h0079e72f_feb79a39,
        64'hffa044df_01d7ccf8,
        64'hffc9d7a8_00d43a0f,
        64'hff348b71_ffe64c8d,
        64'h000e2162_fe67feae,
        64'hff99bd9e_00eea98e,
        64'hffd147f9_ffd2ac41,
        64'hff393439_ffb321f4,
        64'hff516d61_01d14dda,
        64'h00129e16_ffb309a7,
        64'h00a278d6_004693fa,
        64'hfff3e34a_ffef854b,
        64'hff07bb70_0015f8d6,
        64'hff1ea89e_fe00cb7c,
        64'hffe6258d_01d830f8,
        64'hff5aabcd_001ad417,
        64'h007c58ed_01f8a16a,
        64'h0079c2c0_01622084,
        64'h0092cc75_007691c9,
        64'hffc0ccc8_ffda526e,
        64'h001cbe03_01b86677,
        64'h0062602a_ff2516cc,
        64'h00533911_fece221f,
        64'hff20297c_ffbc13e3,
        64'hffb99c94_fef19c7d,
        64'hffe5d3cd_008af30a,
        64'h0079ba37_00bf3991,
        64'hff7e367b_01fcb37d,
        64'h00cade76_ff1163a1,
        64'h00d1b12f_016efdb4,
        64'hff3441f5_fe741497,
        64'h00d3bc99_0076c507,
        64'hff267722_001f2533,
        64'hff908f07_015afd98,
        64'h004dc31b_fe946b7d,
        64'h003364ce_012f92f4,
        64'h008d1439_fef1bc4e,
        64'h00c534a2_01cc2c5e,
        64'h0022bd6e_ff84e4bb,
        64'hffbd07a7_ff77efe1,
        64'h00e76c1f_00520c90,
        64'h00fa2d05_00ec7101,
        64'h00d57957_fec89d29,
        64'h00804b06_00f0922e,
        64'hffa5bd90_fe8e2f25,
        64'hffc1b5a3_0130fa5c,
        64'h00f79170_004f9e7c,
        64'hffcbd90f_fe78c0b2,
        64'h0006e71f_ff62e6dd,
        64'h00617c67_0173d16a,
        64'h00fe5036_ff1b27a1,
        64'h002a9874_fe6f4240,
        64'hff1a5959_0171f2d3,
        64'hffacd2fa_01bc33ac,
        64'h00be4598_ff9347a3,
        64'h00caccb1_015c55b7,
        64'hff4f6b4d_00108828,
        64'hff8685f3_01e6819d,
        64'h00538550_febb52d3,
        64'hffc68b9e_ff1909da,
        64'hff0ad273_014e4f2d,
        64'hff336fc6_0104a339,
        64'h0066e23d_017ed6e9,
        64'h001d82ee_00d195ae,
        64'hffb008c1_00bae5bd,
        64'hff00996c_fe116a48,
        64'h0019099d_019b65cd,
        64'hff549879_fe93eac6,
        64'hff048a57_fe2b87fb,
        64'hff6b998c_ffaf9821,
        64'h005c8375_011bf445,
        64'h005b040b_00ae70aa,
        64'h00cb5425_ff34b3c7,
        64'hff0551ac_011c20c3,
        64'h0090dc6a_014b8c60,
        64'h00d66474_fecf8683,
        64'hff06372b_ffcc2fa4,
        64'hff1d582f_fefa05d6,
        64'hffcdaf4e_0190266b,
        64'hffc693f6_00a9a3da,
        64'h004109b6_fe4f8115,
        64'h001cc778_ff881684,
        64'h005cb375_0196bdd0,
        64'h0066878d_013c0ae3,
        64'hffdd1842_fe989fa0,
        64'hff751b51_fe965407,
        64'hffd6da55_fe071ef1,
        64'hff231d79_0115b64a,
        64'h00bc7cfe_007eeba4,
        64'hff61344c_fe1ecc28,
        64'h000a89bf_fe34e36d,
        64'h0049e85f_fe938696,
        64'hff540293_ffc130ad,
        64'hff32c4ef_01738f72,
        64'hff3ea952_ff9a133a,
        64'hff766cba_feb2e486,
        64'h006e2ac9_007be5e6,
        64'hff427543_feb8f30c,
        64'h00239a3a_01ff62ce,
        64'h005d4b10_00009c08,
        64'hff0be4b5_019b2fb0,
        64'h0022aa9e_01a1d96c,
        64'h00abdaa2_ff66ee7a,
        64'h00b1c27a_fec1c10a,
        64'h00bad355_0189226d,
        64'hff9f2056_fec976f4,
        64'hffa4e5f6_01678a3e,
        64'h001211e4_ff387475,
        64'hfff7ac40_0149c726,
        64'h0021fb60_fe3bc560,
        64'hffd41314_012d49e8,
        64'hffff5e54_01459c37,
        64'hfffca4d9_fe730396,
        64'h009ad133_0191f287,
        64'h00efae7b_ffe1b66e,
        64'hffa1df28_feec7f52,
        64'h00f0ecf1_feadbef3,
        64'hff8675e9_fe6d808a,
        64'h00cc2d84_0134262d,
        64'h00976f2f_fee6d753,
        64'h00aca158_001f7068,
        64'hff748dd1_ff8df61f,
        64'hff219342_00948aee,
        64'hff073b04_0097e7d5,
        64'h00b76fe2_ff29551a,
        64'h00ac8d7b_febae1c4,
        64'h00fe3e77_ff73182d,
        64'h002f24fe_01cb4285,
        64'h00f0c6f8_01b369f2,
        64'hff9eb8b1_0160a7e0,
        64'hffc953fc_ffe5a57a,
        64'h00b1583a_00e49306,
        64'hffbfe104_0119744e,
        64'h00cc2f2a_ff8de743,
        64'h009449f2_fe818b26,
        64'hffcad834_00322379,
        64'hff24c6d3_fff636cd,
        64'hff301ace_014afc6c,
        64'h00b703f5_fed82ef7,
        64'hffd58ae1_fff21c00,
        64'h000be224_ffcc4783,
        64'hff87838e_00f62d6f,
        64'hff2a98a9_fea007e7,
        64'h0072d2d7_fe678f88,
        64'hffa235f9_017ac42e,
        64'hff2d1ecb_fe423c82,
        64'h00264e56_fe7f8ba5,
        64'h00052ae7_fe0e5257,
        64'h005edba0_ff68ab79,
        64'hff3f3235_fe74ead2,
        64'hff8c2417_ff1d7004,
        64'hff1327cc_feb61780,
        64'h008d7a08_002f3f27,
        64'hff4dcd9a_01c91611,
        64'h008e583c_0050e319,
        64'h000ffc7b_ff1499a1,
        64'h00242057_012ca3cb,
        64'hffb4c5fa_0020108f,
        64'hffa10da8_00665c9c,
        64'h0099ae0a_012ab076,
        64'hff8ab39a_017d8e16,
        64'hffbb46df_fe6eb3a5,
        64'hff31c4fa_fe932761,
        64'h00fba98b_007daf79,
        64'hffea3d50_fe004876,
        64'hff6bd65d_005e10a7,
        64'hff806529_01dc2ca1,
        64'hfff5bb6d_0169cf37,
        64'h00e6a4af_fefaa7d7,
        64'h00cf4c1d_007d34e4,
        64'hff34f18e_ffcc171c,
        64'hffd71620_011c1377,
        64'h0096115d_fe547b49,
        64'hff8d5429_ff34a255,
        64'hffbe96e5_01d203de,
        64'hff3119ba_ffd09cb2,
        64'h004a8852_ff019be0,
        64'hff7a4e7f_015986e6,
        64'h000103cf_01945442,
        64'hff3f93d4_fe26d9a1,
        64'hff8cdb5a_007f2ff8,
        64'hff09249a_00a6d653,
        64'hff18d361_fec9f57c,
        64'h008551fb_01a5112a,
        64'h00d0d1eb_0053dd90,
        64'hff9b8d9d_00ef2cb3,
        64'hffe30d75_01d97e38,
        64'hffaa3ee2_01ddbbad,
        64'h00dcf2b5_ffa26092,
        64'hff57c9e1_00e63eb8,
        64'h0003725c_ffe71279,
        64'hff5245aa_00f19415,
        64'h00aa9943_01fa5ce7,
        64'hff33ce28_01fec2db,
        64'h00c1b394_00a1e2b2,
        64'hff284515_019823e5,
        64'hffc5f177_0011d322,
        64'hffdeb5a9_ff3ec4f5,
        64'hffe025be_00e7d32c,
        64'hff45abc9_012e17d2,
        64'hff4d9897_00d14c2c,
        64'h00c6e202_01377ffb,
        64'hff4ad040_ff6d69bd,
        64'h00701b7a_01e55edb,
        64'hff9009cc_ff8e0c3b,
        64'hff0023a0_013f2da7,
        64'h004eb8ce_fff44029,
        64'h00d7b0c8_01e5c0ca,
        64'h004f6678_ff70164c,
        64'h00a41a1c_fe5eecb5,
        64'hff64073e_019205b2,
        64'h000b656c_007681c6,
        64'hff1480db_ff1782fc,
        64'hff83d143_ff882cd4,
        64'hff886034_fe27f9cd,
        64'h00be9487_001c9760,
        64'h007ceb29_01bfd426,
        64'hfffdb64f_ffdab330,
        64'hff9d7d38_fe133817,
        64'h0093aae7_ffffcc5a,
        64'h000946f2_01892bbc,
        64'h00451d7e_ffe186d5,
        64'hffdc2e8f_ff73bd1b,
        64'hffacf3b4_ff9aa271,
        64'hff8c459e_00898506,
        64'hffb398e2_ff03cdd6,
        64'h007a8962_01959826,
        64'h00e660fd_01df0ece,
        64'hff557be7_011c64b3,
        64'hffa2e483_000603d5,
        64'hff9a688d_00830507,
        64'h0098e60e_01692a69,
        64'h006b3cd4_012eeb02,
        64'h0016446e_01f6ef7c,
        64'h00ba12c1_ffa36ec7,
        64'h00c67263_ffa6f40d,
        64'hff8d8f43_fe3dba5b,
        64'hff5444b9_feda6ac8,
        64'hffb1a027_00103803,
        64'h00295f63_0055edae,
        64'h0045ac1a_ff418713,
        64'h00072835_01244a12,
        64'hffd59697_00c73262,
        64'h00e8d1be_ff72f197,
        64'hff0704dd_ff941942,
        64'h004c2334_00716c58,
        64'hffc0c72b_00ad5aed,
        64'hff95bc72_01ceaeb9,
        64'h00730dfd_003441b3,
        64'hfff5d394_fe5cac25,
        64'hfff0d2a9_00fbc004,
        64'hff783b6d_008bb6d9,
        64'h003c12b8_ff62a3c0,
        64'h0098cd3c_00a409ef,
        64'h00bc1c09_fe530f61,
        64'hffd0815c_0105715e,
        64'h00803a44_00595451,
        64'hfffb12d7_010b2fbb,
        64'hffac1a60_fe3feb44,
        64'hff406ada_ffbeca77,
        64'h008bbde7_016f9da4,
        64'hff03e5ba_ff96b59d,
        64'hff4cafd1_018d72f4,
        64'h000b1c30_ff52b68f,
        64'hff8985d5_01da5f3f,
        64'hffd479da_fe7b43f5,
        64'h00108ae9_ff0ff840,
        64'h008cb369_feb4e554,
        64'h0048ae8e_ff6f8450,
        64'hffaf68ed_016e223e,
        64'hff15ce0c_0125e043,
        64'h00944f9e_ff8285b1,
        64'hff7ed72b_ff84b064,
        64'h00740d88_00fe08cd,
        64'h006fa1ff_fec96ca7,
        64'hffd2f8f5_fea85e41,
        64'h00defa18_ff87ea87,
        64'hff06ca37_0153a2dd,
        64'hffed245c_0007ed66,
        64'h0052666b_00b54502,
        64'hff44186e_ff8a23ae,
        64'hff94ca1c_fe63e7e9,
        64'h00bcd16b_ff6c972f,
        64'hff189fa7_00efebd7,
        64'hff4b9558_000a6f11,
        64'h00efe4a3_00f82f4c,
        64'hff6cef86_ffbe4f79,
        64'hff5ba371_017d9b08,
        64'hffd1bd8d_ff6c2601,
        64'hff7d3ab6_01766bfb,
        64'h000d964e_005f8c64,
        64'h0047909f_007f0641,
        64'hffe91cca_ff87ccf2,
        64'h00cbf2aa_fee4687a,
        64'h006d8107_0158d12b,
        64'hff49d2eb_012160fe,
        64'h007d1749_00d86598,
        64'h004e2fcb_fe3305f5,
        64'h003488de_fe87b5f5,
        64'hffbb4261_ffef5aaa,
        64'hfff2148b_fffe0c49,
        64'hff8cbeb7_ffb9e8c5,
        64'hffce7490_ff9179a2,
        64'h00ea9389_001afb6d,
        64'h00270525_01be913f,
        64'h00f556e5_002f9056,
        64'h005ece3a_00bbe140,
        64'hffcc45a0_fe5124ca,
        64'h005565ad_ffae5710,
        64'h003e2250_ff02210c,
        64'h009f2353_ff746ab9,
        64'hffe6a3f5_fe125a3e,
        64'hffd54a2d_fe9879cb,
        64'hffbf1730_01b0b630,
        64'hff3c1ad4_00f3f9cd,
        64'hff8f7a5b_01f1fa16,
        64'hff0b8945_fe0e2bed,
        64'hffe49b74_ff95f84f,
        64'hffa73863_ff779341,
        64'hff63cc4a_fe857edd,
        64'hffb6ed9a_ffef4263,
        64'h00506ffb_01554c7c,
        64'hffb43201_fecbf8a3,
        64'hff8046ab_01fc5459,
        64'h0083a984_00da9629,
        64'hff9ebfd5_ffc3b983,
        64'hfff2d9ee_ff216fa1,
        64'h007f635b_fe9aef5c,
        64'h008126f6_fee58253,
        64'hff412f96_00b52661,
        64'h00736a87_ff753027,
        64'h009be1c6_fea92db2,
        64'h00ff61c2_ff110f67,
        64'hffe9bdfd_fe891d6a,
        64'h009edaed_fece40c3,
        64'hff978a30_009348e0,
        64'h00e1ca81_ff2d6597,
        64'hff521f86_ffd06bb5,
        64'h00b3e294_fe891d5f,
        64'hff06bc33_ff8aaba3,
        64'h0096bdc7_fea744ed,
        64'hff16a783_01069720,
        64'h00dc458a_017bf48d,
        64'hffce4dfa_00814bce,
        64'h008bc658_fe06e55c,
        64'hff4ffef8_ffe8e35b,
        64'h004d7360_ff0c6e74,
        64'hff621161_ff2fceee,
        64'hff7d1810_00898dea,
        64'hffc35d9e_01dbe01b,
        64'h00de64a0_ffb38ea2,
        64'h008706e3_fe0d7766,
        64'hff803246_013b8792,
        64'h004fa401_00a8a768,
        64'h00cc86a5_01a6417f,
        64'hffb5c864_010b1539,
        64'hff6ba211_ffa21daa,
        64'h0064b983_0007444f,
        64'hff5162d1_fee2e51b,
        64'hffe94fcf_ffa46cdf,
        64'h0077aad2_feb46e44,
        64'h00fab3e8_007af071,
        64'hff1f50a6_01171372,
        64'h00aa9579_ffd01083,
        64'hff1622d8_0170b189,
        64'hff335586_fe14806d,
        64'hfffd6ebf_00e3ce08,
        64'h0075582e_fe91c301,
        64'h00bd66f3_ffc86b47,
        64'h0014826d_ff929d5a,
        64'h0057ac29_01d5cc1a,
        64'hff96dd79_007cb622,
        64'hff493f9a_00059829,
        64'h0024ffca_fee58647,
        64'h009a29b5_0179eb20,
        64'h0002e346_001a5247,
        64'hff8853ff_013276bc,
        64'hff0b77ca_0045ab2c,
        64'hfff75cfe_0160725d,
        64'h00251c1e_0042cf44,
        64'h004220e9_fefb7ea1,
        64'h0089b6a3_fecbe788,
        64'h00bf97b0_ff93cba1,
        64'hff7f4540_fe958eba,
        64'h00bd4ab9_013a90e8,
        64'h009c4e22_003747bf,
        64'h0061d1a8_fef5d534,
        64'hffb032c8_ff0d01e2,
        64'hff5412a9_fe923840,
        64'hffb546eb_002b1ee8,
        64'hff3324cc_018c3a16,
        64'hff850bd4_ff7e74c1,
        64'h00e9d09e_fe74e01d,
        64'h004ab8a7_00189f8f,
        64'hff334571_00de19a6,
        64'h00e10cc8_fe40cde3,
        64'h00e628e6_fe61ee6f,
        64'h00be6686_00ac54c7,
        64'hff472bcc_00c6fcde,
        64'hff20e51a_fee923c1,
        64'hffb4e976_fe485c63,
        64'hffae672f_ff2fbe61,
        64'hffa9c8d6_0146f1df,
        64'hff4ec26d_01ddf192,
        64'hff627a88_ffc67851,
        64'hff0b0377_fef6784a,
        64'h0038adf8_014be389,
        64'h00f459cd_ffe24906,
        64'hffa67272_01002c30,
        64'h00aee508_ff1373ba,
        64'hff9ef138_00ecd2ab,
        64'hff018414_01763871,
        64'hffdf1835_fee7e405,
        64'h00e63650_fe5c4c62,
        64'hffea0303_01db9f5e,
        64'h00d65af2_fe10e976,
        64'hff332d77_fe9cad83,
        64'hff323a65_00885455,
        64'hffc0fa6f_00eaf1d3,
        64'hffe9f5b3_ff16dec7,
        64'hfffc5bdb_01e663e9,
        64'h007b0467_feb9f6f6,
        64'hff707a14_00f33da5,
        64'hff4fea6e_fe59bff7,
        64'hff5fd0ce_fe5f32d0,
        64'h00cbb281_005beddb,
        64'h00e200a2_ff630ae6,
        64'h002afe6b_ff01d2da,
        64'hffedb758_01eb772b,
        64'hff2aa45d_feb231cd,
        64'hffbb8018_fef99dc7,
        64'h005ea225_016dc117,
        64'h00307e60_ff9293ae,
        64'hff386bd5_fe71d31b,
        64'h00120b0f_feed35fa,
        64'hff0f1448_ffc68edf,
        64'hffc0bd11_0184bdf9,
        64'h00499310_01911c14,
        64'h002ddaec_01b3fa7e,
        64'h00871f50_01a03787,
        64'hff9b723f_feddae05,
        64'h009abaf5_ff8ede30,
        64'hff8d7224_01a12552,
        64'h007d09ae_ff01b865,
        64'hffe891af_ffe76457,
        64'hff638933_fe924f6a,
        64'hff3e2d02_ffd9a0d6,
        64'h007a4219_ff139cb3,
        64'hffdcd58f_ffc6a75d,
        64'hffe6733f_ff7bba27,
        64'h00059320_0079195b,
        64'h00d1bf8b_fea41990,
        64'h0015651f_01599845,
        64'hffcff3b4_018ee9a0,
        64'h003cafe2_01f49f7f,
        64'hffd5e262_00b9c4af,
        64'h00ee8840_01bd271c,
        64'hff2b0034_01df94be,
        64'h007e8740_01d861e6,
        64'hffa2a2ea_01917e99,
        64'hfff2c0f1_00bf5455,
        64'h0031d0fe_003fbc10,
        64'hffd3a2bb_fe17cea0,
        64'h00649b87_01c6401e,
        64'h001ffa8b_feba5132,
        64'h0074d3d9_008c16d0,
        64'hffe3bbbd_00b02e84,
        64'hff569188_fe6bf9d6,
        64'h00e84380_fe132ce4,
        64'hff90a7be_011ffbd2,
        64'h00ba0c48_ff5dff3c,
        64'h00278a50_01d4bb69,
        64'hffa1526c_ff3f666e,
        64'h0099527f_fe4efe3e,
        64'hff9337b9_ffc55ed6,
        64'h00994f9a_00170f7d,
        64'hffc51175_00c20648,
        64'hff03ff79_017663d0,
        64'h0023d445_00789a8e,
        64'hff751692_00e0f00a,
        64'h00cc3e6d_012667b7,
        64'h00f652ea_ffce362e,
        64'hff18bd62_ffe593fb,
        64'h00c162b5_003d1838,
        64'h00c417a3_00923bc6,
        64'h001061a4_ffecd41a,
        64'h004c3d66_ff47e661,
        64'hff3ec399_ff066222,
        64'hffb978c4_0025969f,
        64'hff6ca12e_00d2d5ad,
        64'h00ef3174_00bd274a,
        64'h0017553c_01a9f3ea,
        64'hffbe0866_0131700b,
        64'h00259d32_feb99109,
        64'hff70ff23_fe99bb13,
        64'hff072989_ff5fce21,
        64'hff905bae_fe5f466e,
        64'hff4f4444_00a86e17,
        64'h000e2dfb_fe483590,
        64'h0071f344_00b48145,
        64'h00cf92f1_fea42fa8,
        64'hfff5d718_0197ab03,
        64'h00d7eb09_00f38f02,
        64'hff5b0224_ff1ede21,
        64'hff4e7ead_fecc72d9,
        64'h0082a2b0_019a7698,
        64'hffb344af_fe182cf4,
        64'h00b6273a_00c21790,
        64'h00f4ef70_0164dfa6,
        64'h007eeabc_ff444142,
        64'hfff95fa9_fee1c537,
        64'h0059c6ca_00cfb833,
        64'hfff8131e_009767ca,
        64'h0004668c_0042fb37,
        64'h00961261_00e48885,
        64'h0092608e_0173b68a,
        64'hff38c85c_fe5e54b7,
        64'h00c76ade_00cfaa98,
        64'h00d3f3dd_00475482,
        64'hffec7c34_fe7fcf80,
        64'h005f9a66_fe914e02,
        64'hffaf6936_019e5b9b,
        64'h00b52f94_011beac7,
        64'h002c93d2_00847ed5,
        64'hff4af764_fecb81b7,
        64'h0029670b_00608f1f,
        64'h00fde2a8_fe1afed7,
        64'h00dac56e_0007cba6,
        64'h00e969f8_ff28af65,
        64'hff744432_004616ac,
        64'hffcf8779_018fc1c6,
        64'h00086cfb_012757e1,
        64'h007f447b_010c84a7,
        64'hff8cb668_01a593f2,
        64'h008d3109_fe7e39e0,
        64'h00ea4e72_ffe84d16,
        64'hff4fcce6_ffd990ae,
        64'hff49e0b1_01759753,
        64'h00e37021_ff705acd,
        64'h001fa751_fed4a28a,
        64'h00a93cb5_00745a3e,
        64'hff4b0738_fe8ba31f,
        64'h00e29d56_01230a93,
        64'h00c3d115_feedcbc2,
        64'hff6cbd3a_0170b1e4,
        64'hffb4f633_ff854a94,
        64'h00016202_01075909,
        64'hff77e95b_01e66fde,
        64'h00e607ce_01e58a50,
        64'hff5e45d5_015cc538,
        64'h00e645bb_ff851803,
        64'hff66bb76_01ecee10,
        64'h005a7ec3_00429954,
        64'hff4197c5_018c9fd2,
        64'h0028ed82_fe3214f3,
        64'hffb97a83_ff498e0f,
        64'hff434646_00727d76,
        64'h00d5501b_fe3126d5,
        64'h006ea045_0060accc,
        64'hff0699ae_fe5d0937,
        64'hff445f0b_fe80ca8c,
        64'hffc67dd8_0102da33,
        64'h005f6ba4_fe9f7374,
        64'hffe6e6ef_ff9dd95e,
        64'hffdb81ce_008b820b,
        64'hff0e82d0_ffa23c67,
        64'hff57d6f3_01b1b35a,
        64'h00ae54fc_fe80528e,
        64'hffba597f_01847aed,
        64'h00feade3_0199402b,
        64'hff3eec04_ff16f5ae,
        64'h004bc05b_01176c6f,
        64'hff124d80_ffdb2579,
        64'hff6c8eb1_fedf8068,
        64'hff7b8c70_ffda6d9c,
        64'h00c2a90a_ffba11a5,
        64'h00ed3782_feff95b4,
        64'h00ca2f3e_00fc73f2,
        64'hff87418d_ffc9bca1,
        64'hffa128d6_ffc84693,
        64'h003c8c79_fe96b3f7,
        64'hff4a1a4a_feff2a72,
        64'hff7f72d0_01446aa1,
        64'hffe25a0c_014ac04b,
        64'h006d6050_0003e3f8,
        64'h00f89515_000e70aa,
        64'hff5c6179_fe61b35c,
        64'hff03fe74_fe5ec55e,
        64'hff7b9fed_ff8d8320,
        64'h00bf3ca9_01f10c19,
        64'hffa0391d_fe20eaeb,
        64'hffbcd83f_ff443e75,
        64'h0095e88a_ff96bb27,
        64'h00f76f0b_fe131c06,
        64'hffab805b_0000a8a0,
        64'hff9594cf_ffe91d61,
        64'hff94a100_004e01b9,
        64'hff8b4d87_fe3231da,
        64'h00b967e4_019a966e,
        64'hff17ce90_0164685d,
        64'hff6b4c71_012588d6,
        64'hffe876ef_fefa3cbe,
        64'hff5e5498_01152b3d,
        64'hff8644f5_01075664,
        64'hfff30b56_fe80d6e3,
        64'h0030a14a_017f357a,
        64'h002bcf08_0094b241,
        64'hffca0dac_ffb62887,
        64'hff8bb2cb_ffaa77a9,
        64'h008114b7_fe697937,
        64'h00c19fd3_00dbc58d,
        64'h0034fd2e_003d7dc7,
        64'h00d9f56e_002b523d,
        64'hff52b431_fee4e616,
        64'hffaaf063_01953989,
        64'h00873552_ff0f64ff,
        64'h00f3b30f_00de8b3f,
        64'hffc129a1_ff60ff17,
        64'h0037b7e8_010b2444,
        64'h00771d81_ffe6655a,
        64'h00129f08_017908b2,
        64'h00981e76_0195a990,
        64'h00638f32_fe76e542,
        64'h00981622_01126622,
        64'hff1b6c18_00903f8b,
        64'hff57aefb_fef95c02,
        64'hfff2264e_fe6736f5,
        64'hffeff443_fe4e8dc6,
        64'hff697baf_0080362e,
        64'hff5bd283_011b32b6,
        64'hff222dc6_01308beb,
        64'hff167978_00ca2d31,
        64'hff006160_0045d73e,
        64'h00fdcf3c_fea5d56e,
        64'hff280634_004e8eee,
        64'h000481c9_01676f0a,
        64'h0095eae0_0072b6c2,
        64'hff918934_ffccb1ed,
        64'hff17abf7_001f4d71,
        64'hff9818fa_ff16e0b8,
        64'hff159aa5_ff9ded0e,
        64'hffd3f17d_fe5d209c,
        64'h00580679_00e55ac1,
        64'h0010c86b_01f49d76,
        64'hffe2637e_016898a5,
        64'hff9e7273_00345ec8,
        64'hffb1cb3b_ff34be8e,
        64'hffbb8afe_ff5dd9d8,
        64'hff6465fb_fe495df3,
        64'hff61ddde_001e9ca6,
        64'h00704af9_ffb7abae,
        64'h0039f4d4_013225c9,
        64'h00642c61_fe9825e8,
        64'h00f6d58d_fefea34c,
        64'hff93db51_015c4b4d,
        64'hfffbf374_fe3d64e4,
        64'h009e3112_ff1895e6,
        64'hff3db2e8_fe851e06,
        64'hff69a35c_0105b52f,
        64'h00e2850d_005cf5d5,
        64'h0046785a_0057f7e1,
        64'h0046f880_fff7f8f5,
        64'hffd752d2_fe97c557,
        64'hffcd082d_fed6ff0e,
        64'hff3e17e3_fe13e104,
        64'hff2b923f_01d7714b,
        64'hffcf7056_ff3216b9,
        64'hffd09610_fe760f06,
        64'hffad0ff4_001cd1fd,
        64'h0042e7da_01932fe3,
        64'h00cd4787_00728a13,
        64'hff2d4036_009e7355,
        64'h0051ab02_fef4b83e,
        64'h007ed0f7_00c49caf,
        64'hff60e115_000dc8d0,
        64'h00291fcc_00e060c8,
        64'hffbc92e8_fff17ced,
        64'hff4c620d_feb0ba78,
        64'h00f0012c_00c4afa3,
        64'h00664bcf_ff9f7b01,
        64'h004da96b_fe78fc24,
        64'h00c72693_fe70c5c8,
        64'hff5c0bd8_fe3dd90e,
        64'h009a632a_fe35126a,
        64'h00d3820c_fe1fa525,
        64'hfffb15fd_00019c34,
        64'h006f0c1d_ff087302,
        64'hffd28bd6_ffffe1cc,
        64'h00b6eb89_004b3eb7,
        64'h005d9c7b_fe005fd0,
        64'h00b487ca_00eaa31b,
        64'h0096abeb_fe007457,
        64'hffc9c436_01462495,
        64'h0029ce01_fe7f639d,
        64'h0087fa9d_ff5414d8,
        64'hffe8aad4_fe37b4d9,
        64'h0034d40a_fe0cd19c,
        64'h002462c7_0161dc94,
        64'hff69d633_fe390c5f,
        64'h0052704b_fed9e879,
        64'hffef990f_ffc609e3,
        64'hffe72579_00cf56e0,
        64'hff5b7dbf_fe9e74e0,
        64'hffc710f1_00f5ba3c,
        64'h00f2f2ca_ff00e985,
        64'hffa47b01_00ea09f0,
        64'hff67b518_011452c0,
        64'hffa4669d_00ef4fc0,
        64'h00bbe717_fe5ba384,
        64'h00003c82_00326916,
        64'h001f4ec8_00fd8933,
        64'hff96b225_ff17b784,
        64'hffbd2f56_fe7ae7a9,
        64'hff19f480_01bf8dd3,
        64'hff0ce532_00fbfdbd,
        64'h00e5da2e_0052304a,
        64'hffbc8bd9_febdb5eb,
        64'h00ef86bc_ff5195ba,
        64'h003aca30_ff671929,
        64'hff9c8716_fe0aa885,
        64'h004811b8_00e2377b,
        64'h0078e3fa_01a0c15c,
        64'h00a15142_009ae7bc,
        64'h0077bf1b_fed32b58,
        64'h00f4c534_00bfebcc,
        64'hff373293_fe3dcbad,
        64'hff515462_00354ce4,
        64'hfffabcc0_00f42772,
        64'hffe0379d_feec8d3e,
        64'hffd2ff33_ff3e817f,
        64'hffe6949e_0121ee60,
        64'hff0d10d6_fe523c68,
        64'h00048f7f_01b7b2ad,
        64'hff795015_ff68a362,
        64'h006e4e88_ffd30fd8,
        64'h005b6d8d_0026cfa1,
        64'h00093c11_01e0f6d0,
        64'hff48b650_fecebdfb,
        64'hffbe2b7b_016ca37a,
        64'hff87de86_010bed3a,
        64'hff395d6f_01f78f84,
        64'h00739fa0_fec80312,
        64'h00c2c250_fe4b193b,
        64'h0038d0e6_00f4a064,
        64'h0009488d_ff3bc2af,
        64'h00503b47_019a2109,
        64'hffd4d441_fff9b7ca,
        64'h0044f155_01112c4c,
        64'hffdfc441_00c47b4f,
        64'hff579341_011bddfa,
        64'h00191e33_00dde59d,
        64'h00e834a7_ff2b6aeb,
        64'h00ff01d1_01712192,
        64'hffc2c815_015cb735,
        64'hff36f5a0_ff9ed690,
        64'hff9ebdfd_016e5968,
        64'hff2efcfa_fe57cfb2,
        64'h00ce418c_ff08b351,
        64'hff79c8d9_01c7bee1,
        64'hff27db52_011a5be2,
        64'hffed4c62_0087e5c3,
        64'h00dccdaa_fe081bee,
        64'h005fb709_01b2d808,
        64'hff703bf8_fe4bc754,
        64'h00ac546f_fe82976e,
        64'hff4a8632_ff21aed6,
        64'hff645061_ff418a4a,
        64'hff0a6706_00d09380,
        64'h0053ca69_01383922,
        64'h0006f4a1_ff38402d,
        64'hfff7193e_ff7eb9ec,
        64'h008ff749_fe89aeb1,
        64'hff75098f_fef77a3c,
        64'hff8b5488_01b7f946,
        64'h00f1e3b0_0172e328,
        64'hff9360ab_ffcdd83a,
        64'h00ead64c_fe28539e,
        64'h00a26e6f_ffa54401,
        64'h00c26b32_fe75a02c,
        64'h00cc2390_00fb9c3a,
        64'hff486d0c_00866908,
        64'hff34105d_014232c1,
        64'hff55704e_ff48042f,
        64'hff12b8cd_004c5436,
        64'hff76659d_01ef8f75,
        64'h0092396e_ffb00bf0,
        64'hff193316_01860a28,
        64'h00201784_ff75ae30,
        64'h003abec1_ff790e52,
        64'h002f3580_01a4e931,
        64'hffa16eb8_0149e3c3,
        64'h00e3084a_fefcb4db,
        64'h00c22358_fef8790b,
        64'hff61afe8_ff1a1960,
        64'hffeaed3b_01de9e46,
        64'h0082b755_0161c4a9,
        64'hff500692_fea49e39,
        64'hff85c28c_0046e672,
        64'hff14dc6c_007001e9,
        64'hff66c64b_fe196809,
        64'hff82b0bd_01c74c21,
        64'h003b8469_fe603de8,
        64'h004a449a_fe99b2f6,
        64'hffa8879b_00d4fd5f,
        64'hff37d7ab_016c7c1b,
        64'h00263811_019cc075,
        64'h008ccd0a_ff580710,
        64'hff8fc1bb_01a6e146,
        64'h00d9a6d9_016e44d1,
        64'h00869ee0_014bea52,
        64'h00bca47f_ff3f3ae0,
        64'h00a9a86f_fe1891ec,
        64'h00c073dc_00a13d11,
        64'hff0f8dec_fe2d5d1c,
        64'h00e1936a_018144be,
        64'h002dec33_fed70f2c,
        64'h00073619_000c93d3,
        64'hff8a34e8_00a643cc,
        64'hff697e22_ffe83675,
        64'hff69607a_fe3010ff,
        64'h00b25960_0076b1be,
        64'hff99088d_ffd37a82,
        64'hffc654f1_ffb5da89,
        64'hff18456b_ffa1d4dc,
        64'h0016699a_00f5a82e,
        64'h00dfa8cc_fe89927d,
        64'hff8557ed_013d1def,
        64'h0008050e_005675b9,
        64'hfff682e4_ff68d7e8,
        64'hffb574fd_01f9df4b,
        64'hffdbd7c7_fe5e8174,
        64'hffa0d9c5_0086d4ce,
        64'hff732772_000c1ad3,
        64'hff9ce5a2_ffe73272,
        64'hff237678_ff1461c9,
        64'hff5dc6e2_ff548510,
        64'hffee52b2_fe532d92,
        64'h00359213_fe4732d3,
        64'hffa23f97_ff8f626f,
        64'h00dbafbc_fe8c2bcc,
        64'h005e128f_018adbb4,
        64'h0088bd51_fe34cccd,
        64'h004d175d_017983e9,
        64'hfff73e11_ffce405f,
        64'h000e84d3_00ed89df,
        64'h00c89af4_fed7e7c6,
        64'hff0d1c1d_fe545b16,
        64'hff264a65_003c6ff7,
        64'hff1620c0_fe1534d7,
        64'hffa7cef9_ff2b4f29,
        64'h000de052_01f47944,
        64'hff5d6754_ff31f467,
        64'hff13ab47_ffe8f7e9,
        64'h00a3e1f2_00165f39,
        64'hff94caf8_002ed8eb,
        64'h00f994b8_fe1e6f8f,
        64'h006862d1_00983678,
        64'hff5f9691_fe066215,
        64'h007e642d_0177a5a7,
        64'hffbbc92f_016139b7,
        64'h00e97790_ff887ebf,
        64'h00b975ed_ff3f5f75,
        64'hff3578b5_014e0583,
        64'h005b61e9_0011a212,
        64'h00429706_fe35a053,
        64'h00c1c970_ff977787,
        64'hffe438d6_0100ecd5,
        64'hffa934e5_fe52d159,
        64'hff975e54_01b3a3b4,
        64'hff062fff_008472de,
        64'h00f9defd_fe0a2daa,
        64'hfffff4f1_fe1f0027,
        64'hff0db0fc_fef7e404,
        64'hff1e2ad5_fed39d1f,
        64'h005e9b8e_fe168643,
        64'h004525e6_fe129431,
        64'h00214cef_ffdb2efd,
        64'h0054f63d_01e08194,
        64'h0079e72d_ff58188f,
        64'h00ebaa50_ff4d690a,
        64'hffde6f34_febfab44,
        64'h003fb6e9_fe37de4c,
        64'h004bd71c_ff136c7c,
        64'h00fd0583_fe8c1b84,
        64'h00d4c4d8_ff884fd6,
        64'hff570e90_fe6fb74c,
        64'hffe82836_fede4718,
        64'h00f3d675_011fc8c0,
        64'h00a2efd2_004b613f,
        64'h00c2c90a_01f3fe19,
        64'hff838a8e_00ea33ef,
        64'hffb838ab_fffb9c2e,
        64'h001ce8fb_fe86cf9d,
        64'hffd9589e_00950efa,
        64'hff03f4f2_ff37d29c,
        64'hff3e41ff_019a6313,
        64'hffaf63c1_00aff431,
        64'h0097e08d_ffd48975,
        64'h00c10d11_ffb411dc,
        64'hff194ec2_ffa7a956,
        64'hff8c3850_019689bc,
        64'h00ed908b_ffe2d887,
        64'hff5468f3_ffa8b8ee,
        64'hff61688a_ff7d8784,
        64'h00bba848_ff836583,
        64'h0022702c_fefcfbc6,
        64'hffb849aa_ffe3300b,
        64'h00c252e8_01d6e347,
        64'hffcc1523_ff35ae89,
        64'hffebf7f7_0134e6dd,
        64'h00ae5f1e_00680800,
        64'h00c65c93_01abbc55,
        64'h00f57a5e_012c8891,
        64'h00b75709_01a200fd,
        64'hff59d334_006ee83a,
        64'hffcb9b84_fea62d38,
        64'hff5b09c9_ff5db434,
        64'h00349ef9_00d87bb9,
        64'h00386fda_fec6adbb,
        64'hff8bc176_ff526374,
        64'h001eab29_003cae1f,
        64'h00fa07ae_005ab4e4,
        64'h004e826c_fe32d1cb,
        64'h00fb0aad_0190288c,
        64'h00f45b9a_014dc26f,
        64'hff623a3c_011f330b,
        64'h0026ff10_00bf932e,
        64'h009db192_012b0c3d,
        64'hff5e3b76_ff4f63c1,
        64'h007b4aa1_00de7499,
        64'h00064626_fe40898a,
        64'h00f95dcb_0076816e,
        64'hff9545ff_01181bc1,
        64'h000f24d7_fefc4b03,
        64'h001fac7d_fe8bbe71,
        64'hff9393b3_012ea9bf,
        64'hff3daff2_ffc1050c,
        64'hff542468_01d0da4e,
        64'hff5c8626_fed248e5,
        64'hff3f8800_000a261d,
        64'h00e20161_00c10909,
        64'h00c0ee8c_fe142557,
        64'hffd9a295_fff6ed7d,
        64'h00b37f80_fecd5d05,
        64'h0000c474_000a9ff5,
        64'hffa4f2b1_01ddcb2a,
        64'hffdba160_0108773d,
        64'hff2677be_fe267ff6,
        64'hff2895c2_ffa203b9,
        64'h00462a3c_016c011f,
        64'hffd73dc3_00a7366f,
        64'h001831b1_00b41ba9,
        64'h00673588_fff38653,
        64'h00588d06_011336d4,
        64'hff7b6841_00673f75,
        64'hff960395_ffc74686,
        64'h00bb117a_ff46f6c2,
        64'hffc9b91f_01abe671,
        64'hff66cdf0_ff5c2f66,
        64'hff07f808_0023b4dc,
        64'hffeb2c45_fe18d5f2,
        64'h005beae4_ff56907e,
        64'hff6f4a2b_00f6ae56,
        64'hff2342b4_ffa57cde,
        64'h00447613_014aac23,
        64'hff0bf945_fe5c3b4f,
        64'h00eb68ed_ff61766f,
        64'hffb0a031_00e6bad9,
        64'hffec11c5_01f91254,
        64'hff64d120_00220d10,
        64'h0090a9d7_0052acd5,
        64'hff7d0f53_fe295ac0,
        64'h0098d121_018f7b2c,
        64'hff566592_00b1ea92,
        64'hff36b788_fecbb08f,
        64'h00f9bf84_fe17752d,
        64'h009360b7_00b4d67d,
        64'h00410437_fe66feb2,
        64'hff0c7cb2_fff665f8,
        64'h0016aa6d_fec79399,
        64'h00e45de1_01ca0318,
        64'hffdf17c0_00aa48fb,
        64'h005d6e69_ff700dfb,
        64'hff8c7abd_0026bae7,
        64'h00ad1910_fe68d25d,
        64'h00ba9245_fee29253,
        64'h005bd2b2_fef9dd37,
        64'hffa510e4_003e9144,
        64'h005b03d1_fe9a256e,
        64'hff94f656_fe7e697a,
        64'hff05e746_002be191,
        64'hff8199fc_fee6aa81,
        64'hff9271b1_01e41e16,
        64'h00f30d57_00cb90a7,
        64'h003c5480_ff5b7376,
        64'h00f6a56f_001cad3e,
        64'hffd82d0a_ff5971a6,
        64'hff323431_0022cfe8,
        64'h00cfeb55_feb2368a,
        64'h000cdf03_ff34d9c2,
        64'h00e72b92_ffa4af3b,
        64'hffc7eec8_fed06002,
        64'h0081d4ec_ffbd232e,
        64'h00eb1236_0116e835,
        64'h00fc2f5c_01c59c13,
        64'h008e4d71_0175038e,
        64'h00726eb0_01ba47fc,
        64'hffe81b10_ffc66c0c,
        64'hff8f6623_fe2d2851,
        64'h0004c235_006ebfcd,
        64'h007966ae_ff06fdc9,
        64'h00e2c296_ffad42cb,
        64'hff87da5b_fe0aa76f,
        64'h0000046d_004a31c0,
        64'hffbc6025_00009e02,
        64'hff0321cb_00a4ca7f,
        64'hff6c28da_fe901743,
        64'hffa4cc50_fed081dc,
        64'h00347e37_ffcf8eee,
        64'hff7eb979_006feca8,
        64'hff463c29_fe359cda,
        64'h00f2bf02_fe06b720,
        64'h001ae90a_fef4136f,
        64'h0074ea42_ffddec5b,
        64'hff6ea624_ff176ea2,
        64'hffec6958_fe7fdbe3,
        64'hffd177b9_01d31076,
        64'hff276b5d_ff7213a0,
        64'hfffc2f20_010d514e,
        64'hffdc9358_ff275d3b,
        64'hffe8985e_ff3596f4,
        64'hff85522c_016d6557,
        64'h00fd9392_0070cb20,
        64'hff99b829_01d8fb46,
        64'h00e9413b_018bee9d,
        64'h00e94d49_fff4d878,
        64'hffa1e30a_ff35b893,
        64'hff190eb1_008c85b6,
        64'hff854958_0138aecf,
        64'hffd6a910_016a3f40,
        64'hff2fab8a_ffc4c301,
        64'h008e0fe6_ff45bfd5,
        64'hffbfb7f6_014b710c,
        64'h0039f38b_ff0cdf06,
        64'h00d43419_015a11f1,
        64'h00e36ee4_0124a509,
        64'h00a48c50_fe530c4b,
        64'h0032c342_ff8975f5,
        64'hff08d6b6_ff601744,
        64'hff2ad2a4_fea22225,
        64'h00e12bd3_ff7494ba,
        64'hff303215_fe0dcf18,
        64'h008dcf1a_015c6920,
        64'h000efb72_fe61bf5d,
        64'hff574137_01ffe6c8,
        64'hff2d82dc_fe0898d9,
        64'h00a73d1c_00ca0db6,
        64'hff92946a_ff7cfa9b,
        64'hffedfb30_019da60d,
        64'h00da0c8d_ff7c7cc9,
        64'h0002932e_ff65015e,
        64'h00f37e35_fe0bee6a,
        64'hff635ec4_006058bf,
        64'h00d965f5_fe5ea5c0,
        64'h0027b6e5_ff896d17,
        64'hfff7afa9_0008ea2c,
        64'hff72bc3e_00d21d63,
        64'h002e6ae0_ff5745c6,
        64'h00fdaf5d_fe5da4ea,
        64'h0025b304_ff9baefb,
        64'hff504234_01eb2181,
        64'hff496000_ffe0d457,
        64'hff36b82d_01511c9a,
        64'h0040bdcf_fffde043,
        64'h00834054_00f7ba73,
        64'h0001a94f_00ad2d08,
        64'h009236e6_0092595e,
        64'hff9e4981_ff589e05,
        64'h008ef084_003aa73f,
        64'hff6e7ff6_fee26728,
        64'h0072ef06_fe656a28,
        64'hffd7c923_ff69d025,
        64'h00a81059_fe70220d,
        64'h0011cf4c_008a763a,
        64'hff79e53d_ff646cfb,
        64'h00e7a57e_001a1a1c,
        64'hffc639a6_002aa810,
        64'h00bea32d_01c7db77,
        64'hffae241a_01b20a7b,
        64'hff3ee90a_001aef18,
        64'hff64d8e5_00d01742,
        64'hffe371c2_ff002ac8,
        64'hff664aa6_015b4841,
        64'h00ccff1e_fec7a40e,
        64'h00a5a8c1_fea348cb,
        64'hff51d3b2_ff854ff0,
        64'h004981a6_ff85bc9b,
        64'h00d757a8_ff034a97,
        64'hff49eee5_00a6ced4,
        64'hff536514_ff141188,
        64'h0097bcd4_fe22ff82,
        64'hffbdc15d_fed5facb,
        64'h005c4fb2_ff7483dc,
        64'h004868c2_ff710aa2,
        64'h0096d508_fe3c6772,
        64'h00a32c89_001f893b,
        64'hffe3ba70_fff57623,
        64'h00489f31_fe8d5bb6,
        64'hff33db88_018647c3,
        64'hffbdab30_0179d109,
        64'hff55af77_ff6dd07c,
        64'h0030be85_00c6a5b7,
        64'hffe4dffe_fff927d5,
        64'h0015770e_01b6dea2,
        64'hff426c1d_003074d4,
        64'h00cda6ab_00be7af3,
        64'hff62d1ae_ff8779e7,
        64'hff86b34f_001c793a,
        64'h00a82995_ff14ef9d,
        64'hff4eaaa8_fe724a13,
        64'hff3c1122_00b06cf6,
        64'h00886752_ffd24fb6,
        64'hff14c66c_fe234992,
        64'h00c664eb_0192e639,
        64'hffc99185_00ccd72a,
        64'hfffbd9c7_ff61483d,
        64'hffcc4d6f_ff81ec4d,
        64'hffd2ef16_ff81302e,
        64'h00650bbb_004a144b,
        64'hffb91012_0124cf79,
        64'hffa49467_fe2f34ec,
        64'h00e6df5f_015aee39,
        64'h00110f4d_015299fe,
        64'hff3dfa72_015905f4,
        64'hff7b7803_0196b25a,
        64'hff360435_fe6a6b4a,
        64'h00a5626a_01f501fb,
        64'hff2b0837_008f7824,
        64'hffe6d6e0_01a65ca4,
        64'hff4030e6_0170f839,
        64'hff14759c_fe5e7de2,
        64'h00467e09_ffe2231e,
        64'h0036f5eb_01d1d52b,
        64'hff65cba8_0051590a,
        64'h00c27d94_fed31b8a,
        64'h00254aaf_fed0afac,
        64'h00cf404c_00b83eb9,
        64'hffc5af39_fe2e8411,
        64'h004d54a7_ff623b0e,
        64'h00d55bee_013a883d,
        64'h00f66569_0150f43f,
        64'hff464ffa_012a4dd3,
        64'hff824cfb_ff61f2b2,
        64'h00680364_01b17bf4,
        64'hffc06bd6_0075cba5,
        64'h00130d60_01f623ab,
        64'hffa5a0da_000f11bb,
        64'h00fdaa95_ff44a32e,
        64'hffd5a16b_ffe5ba44,
        64'hffac9076_fe1a246a,
        64'h0025904c_fff38119,
        64'hff538cb2_fe26cc22,
        64'h005f9126_005bfb96,
        64'hff2b9865_ff87d8ab,
        64'h00b7610f_013b32ce,
        64'h00832487_01812204,
        64'h00f612fb_ff3666e1,
        64'h0006ef3f_fe79dba2,
        64'h0085deff_fe36dcb7,
        64'h002763b7_01eaa592,
        64'hffa8be85_ff895fc7,
        64'h00e47468_fe8a1528,
        64'h000aafcc_014f7fa1,
        64'hff70702c_fef32123,
        64'hff3be96b_00a7bdda,
        64'hff0e9959_feac4d91,
        64'h00b3b310_01c619d4,
        64'hff537763_fe7fe3f7,
        64'hff16d1b1_011361cc,
        64'hff4e57f1_ff931d82,
        64'hff578a24_ffa7707c,
        64'hff612550_fec82a8a,
        64'h00eff595_ffda8e7a,
        64'h0043974f_ff76f1cb,
        64'hffc995d9_ffde5c61,
        64'h0068fa87_ffb58bc2,
        64'h008d0c32_ffbb2f02,
        64'h00f068af_00a4283d,
        64'h003b717d_01eb426d,
        64'h000c0bc3_00b36a3c,
        64'h007af6e8_001386fd,
        64'hff4d25eb_015265b8,
        64'hff1bedb9_00e0f177,
        64'h00c0b64b_01205392,
        64'h006db101_00561855,
        64'hfff6653c_0140d4bc,
        64'hffe75a0e_fe171fdc,
        64'h00ed4898_00c5d975,
        64'h00d53be2_ffd07ef5,
        64'hffed1368_009fe0a6,
        64'hff4eaccc_fe912b77,
        64'h00a29652_fec8fec3,
        64'h005f108c_fe9879a2,
        64'hff3b6092_ff9d167e,
        64'hfff2ac48_003405c4,
        64'hff3848a8_007665cf,
        64'h009ba270_ffd2dbd4,
        64'h00a3f12c_fe51b987,
        64'h0049f056_00bf0fa2,
        64'hffd7de5b_ff7e8005,
        64'hffeefe1c_01d17b78,
        64'h00ce198e_01fb2de2,
        64'hff03f14d_ff6e249d,
        64'hff41443f_00104f51,
        64'hff327507_00bf6926,
        64'hff0c4704_015172e3,
        64'hff09232c_00e96ff2,
        64'h0043f320_fed9b011,
        64'h002b4f8b_0134cdee,
        64'hff87bab0_fe1f45e6,
        64'hfff8eaf7_01d2e48f,
        64'h001eba15_ff34815b,
        64'h00dfcd58_ff17c824,
        64'h00fe078e_00b8f70d,
        64'h000ea902_00fbf685,
        64'hff91d03e_0093f1cb,
        64'hffa6c55f_00266512,
        64'hff8665cd_ffb60962,
        64'h002b8cd0_ff685277,
        64'h006a95e0_00b48a48,
        64'hff42b477_0191cb72,
        64'hff7ae681_ffb7510b,
        64'hffd55b3b_000cd994,
        64'h005bee1a_01c03dd3,
        64'h0027c811_019f5168,
        64'h00fcc747_ffc79aba,
        64'hffa01b4a_feda7c1f,
        64'h005045c8_fe782522,
        64'hffad75db_00bea46c,
        64'hff669f41_008f8eed,
        64'hff1ef6d9_00866889,
        64'h00707dcd_00493df5,
        64'hff22a177_01e50dad,
        64'hff253887_fe2e147b,
        64'hfff949df_0123b81e,
        64'h00c51ca0_ff127de7,
        64'h000867f8_ff737174,
        64'h0040030c_ff41c6d8,
        64'h000aae5a_000ee8d4,
        64'hff6488a5_feab3d24,
        64'hff869c04_fe367825,
        64'h000403c5_01f3dce5,
        64'h00753ae9_ffd944be,
        64'hffbd6a6a_ff322aca,
        64'h00a3bd2a_00d4d18c,
        64'hff1798d7_00436c61,
        64'hff297a88_fe6fa0fe,
        64'h0035fac1_00e82972,
        64'h00b0ef32_ff146ea8,
        64'hffd399eb_fe180160,
        64'h00ef768b_000498a4,
        64'h002dfd2b_005dda61,
        64'hffcb6ab2_0087ba0b,
        64'hfff1a6f4_ff761775,
        64'h00ba735f_feb10d90,
        64'h009d5f36_00359654,
        64'h00384d8b_fe283982,
        64'hff0d5488_00e14444,
        64'h001c69f4_00ace183,
        64'h008d8e2b_ff6721c5,
        64'hffa45d48_fec2d3db,
        64'hff06a9d4_0046a5d6,
        64'h00f5a857_ff7d2919,
        64'h0029380e_ff3d784e,
        64'hff368257_fea09b7b,
        64'hff90bd34_ff04d9c3,
        64'h00a5c8fd_011b1067,
        64'hff348e69_ffb513e8,
        64'hff92a6c1_0031c06d,
        64'h00de0798_ffccaabf,
        64'hffed5be7_00209e25,
        64'h00700286_011bcd54,
        64'hff07fc1a_00f587cd,
        64'hfffde609_fff9c30e,
        64'hffa5d94e_00229a59,
        64'h0001bb49_015eccdc,
        64'h00ee7263_006b383c,
        64'hffc6316a_0107e3ec,
        64'hfffbdc80_016758cc,
        64'h0025f8dc_0046fc78,
        64'hff2079b2_ff243e6d,
        64'hff8a5d83_fe6ab0b3,
        64'hff999962_007dd9d6,
        64'h00113ee0_01d82d51,
        64'hff5321e6_ff6c0290,
        64'hff237d3e_00d5db1a,
        64'h00caf278_ffb28b4f,
        64'h000a970a_ff3e9718,
        64'hfff710f9_ff5dc2aa,
        64'h007c39ef_fe84d437,
        64'h00e2eed2_ffce4d96,
        64'h00692787_0188fee3,
        64'h00ae10c3_fe20e114,
        64'h00bc6de4_ffab143b,
        64'hff14dc31_feecab75,
        64'hff80718b_fee7bc8c,
        64'hffdd5f82_003488c7,
        64'hffe5d3a3_0058aedc,
        64'hff5e5a0a_010bb3a0,
        64'h0012be1f_fe96e3a3,
        64'h00d5dd26_ff4fe4e3,
        64'hff6c44ad_fed712de,
        64'hffaffecc_005b2f64,
        64'h00bbd45e_0085ba83,
        64'hff0b26d8_fedb7470,
        64'hff179bad_ff57923d,
        64'h00e7e3c2_ff41424e,
        64'hff49e45e_01154557,
        64'h00f450f1_01112781,
        64'hff37f999_01f37446,
        64'hffa07038_fee15deb,
        64'h00622d7d_00170b9d,
        64'hff89668f_ff24b8a2,
        64'h00db44ad_01dec068,
        64'hfff9e2e4_0092428e,
        64'h00063578_00463218,
        64'h00c93773_fefe5eb9,
        64'h001858bc_01cf795f,
        64'h000a93b0_01921e1a,
        64'h003b61f8_ff02210a,
        64'hff443b1b_fe0758b2,
        64'hfffb0dae_016d67ad,
        64'hffbf0fb9_fe096363,
        64'hff97a9d5_fff10177,
        64'h001738e9_001191e6,
        64'h0084ff8b_01f8b5e1,
        64'hff34655b_fe6b400a,
        64'hff0d8c38_01f94838,
        64'h0036cfa0_fe00cbfc,
        64'hffab6576_fe7a0964,
        64'h00cfb850_0095fecc,
        64'hffe24805_01100dad,
        64'h005cd15b_009abf9e,
        64'hff4c352a_002eb079,
        64'hff533828_fe998dc2,
        64'h00777064_feac9ef0,
        64'h000ef990_018f5870,
        64'h00ea0866_011a73d0,
        64'h0023cce3_010c85ee,
        64'h00959581_015fa966,
        64'hfff8d948_ff8f57e3,
        64'h0063f0b7_ff73131f,
        64'hff6c4f72_ffea32a7,
        64'hff33dae3_ff0b7019,
        64'hff6cf047_fe51bc90,
        64'hff7b7ba5_ffb488b3,
        64'hff7b3f11_01096ebe,
        64'h0012a3b4_00da64b4,
        64'hff246d9b_01ec0dd0,
        64'hffed5787_01e99de9,
        64'hff7f4d6a_feba4793,
        64'hffbe9300_ffbd5e4e,
        64'hff8ca9d9_ffee1a41,
        64'hff07538f_0028a06d,
        64'h00e9704f_00047f37,
        64'h008caf3f_fed711a1,
        64'hffaaec41_fe1e43fd,
        64'h00243d7f_0106c119,
        64'hff5264a3_fe7324f4,
        64'h0050165c_00326f32,
        64'h0092f845_ff4bdc5a,
        64'h0071b1b9_01d487fa,
        64'hffe8557f_01f30b98,
        64'h00933825_ff0542ca,
        64'h008c7224_00bba2a5,
        64'hfff11a5f_0118c14c,
        64'h002d2467_01d0655e,
        64'hff5182bc_01cad202,
        64'hff58c77b_01dae8f1,
        64'h0079b303_001ed10a,
        64'hff0fb545_0067f22d,
        64'hfff67f84_ff4c081e,
        64'h000c6f0f_005d62b7,
        64'hff3aa2d0_0038df28,
        64'h00483946_fecaafb0,
        64'hff7a9fe3_ffc2f20f,
        64'hff6d3224_012df38d,
        64'h0023ada8_fecc01d2,
        64'h00ef2835_fe895ca6,
        64'hffbfc1ce_fefa80b3,
        64'hff9932ec_01571c44,
        64'h0068b01a_0195d792,
        64'h0006702c_feb9a02e,
        64'h002a4851_fe02c09a,
        64'hff0d0d2d_fe8c3fc8,
        64'hff499a77_006f6f9e,
        64'h00778662_01b39c0b,
        64'h005346bd_fe1233b3,
        64'hff185421_00351c59,
        64'hff3b2b92_fef39339,
        64'h00fa412c_fe8255c9,
        64'hff4b3326_ff79f397,
        64'hff25c79a_00b84763,
        64'h00c343f8_fed2e513,
        64'h000fcd1a_febc182d,
        64'hff2c633a_fe56a355,
        64'h00ae480f_01bedefd,
        64'hff910e57_013d800b,
        64'h00c20181_ff526e16,
        64'h004cc7fc_01af0a50,
        64'h004d088e_004638ca,
        64'h0098fd5b_0157c81a,
        64'h002b545c_ff166f23,
        64'hfffce9a8_01a8d838,
        64'hff62618f_002fa34b,
        64'h0043bf27_00eea82e,
        64'h00813c68_0088e8e5,
        64'h00ebd8a8_fe5b0366,
        64'h001b8734_013b19ea,
        64'h00633cde_fe93c765,
        64'hff673ae0_01635961,
        64'hff76a1c9_ff18256a,
        64'h0003c7c0_fe5872df,
        64'hff7623f0_ff95a3db,
        64'h00f24a61_00094db9,
        64'hffd6fbaa_ff9ee2eb,
        64'h002c3624_018e025e,
        64'h0001c6ca_ff6d01dc,
        64'h005cef67_01dc9a1e,
        64'hffe59b7d_ff1d01a5,
        64'h0058a208_fe01acc9,
        64'h009add43_ff6dc168,
        64'h0023679d_ff54b610,
        64'hff2baf31_00547e9e,
        64'hff319b4e_fe844972,
        64'hffac623b_00e62df2,
        64'hffa9594c_0186f50e,
        64'hfff9551a_ffd9ca94,
        64'hffd357cc_017f3173,
        64'hff749c6d_fe2ffcfc,
        64'hff01da5b_ffdb6d0e,
        64'hffc8507d_00968ca6,
        64'h00f30a35_ff78df93,
        64'h0070ccd9_fe1262b3,
        64'hff67a28b_ff8ff520,
        64'hff49f086_ff5dfe57,
        64'h0078b583_00beb9a6,
        64'hff6d76ac_01f75ef5,
        64'hffc758af_01d465e2,
        64'hff8d5452_01d54d52,
        64'h00b22574_ff56a04f,
        64'h00fb1db0_ffdfb84e,
        64'hffbb2d61_ff693348,
        64'h00d2e2a1_0004d5ce,
        64'h0090b283_0022bd18,
        64'h00a7cf6a_012e2725,
        64'hff53c8ac_fe0ec552,
        64'h009e54fc_fff70cb2,
        64'hffae989c_01803a7d,
        64'h00fb8a43_ff1b63bc,
        64'hff38ae70_00feac1f,
        64'hffa05e7c_ff3ed06f,
        64'h009cba83_fe2165f1,
        64'h00a62e34_fe8aef26,
        64'hfffe71a2_ff0efdf0,
        64'hff34b4e9_00683aa3,
        64'hffac8dc8_01ec4caf,
        64'h00b6a16a_01907c5a,
        64'h00e9ab89_009d806b,
        64'hff5f3345_016610c1,
        64'h00300f67_016c7fd3,
        64'hff4c7471_fe640193,
        64'hff29d32d_010f9e56,
        64'h0076018c_fe9e7614,
        64'h00aa99d8_ffc486bb,
        64'hff835de1_fff3f8fc,
        64'hff854e5f_fefbc5c2,
        64'h00ab9114_ff54a701,
        64'h00be63dc_01258593,
        64'hffba2260_00a4c59a,
        64'hff69a705_00e93c39,
        64'hff5dc46e_019cb6df,
        64'h00c98573_000a9f26,
        64'h0052d189_feb39075,
        64'h006c9718_01d51b9f,
        64'h00e34c9f_01531a53,
        64'h00cce357_ff900e57,
        64'hff0f5b2e_009b75fe,
        64'hff6c7533_ffc434d4,
        64'hff58b868_01e42bf6,
        64'h00c970d0_00adbb36,
        64'hff8efab9_ff21bc51,
        64'hffa670a6_ff89ef25,
        64'hff33edf6_ffb304b8,
        64'h00ef7563_fff512f9,
        64'hfffb11ca_feef1191,
        64'hff387304_ff93f0d4,
        64'h003de819_007877f2,
        64'h000aab31_00615314,
        64'hff0ef52a_01266e52,
        64'hffe1b075_ff23caac,
        64'hffcee3e5_008d8ef3,
        64'h000d3e28_fed8dbbc,
        64'hff14b3f8_00a5602c,
        64'h00a195b9_0070c557,
        64'h00c75997_00b16272,
        64'h00ec7092_0176dd26,
        64'h007bd67c_0042cc9c,
        64'h0008314a_fea758f3,
        64'h00d97de9_feb9402b,
        64'hff93eb3d_00a20eae,
        64'hffcafe4c_00a47034,
        64'hffb50ceb_002d9068,
        64'h008e6d5d_fea7f133,
        64'hffb5c41d_01721fcc,
        64'hff5f3020_00e73bea,
        64'h00896f4b_012d47cc,
        64'hff042762_01150951,
        64'hff7fc647_0156f9a2,
        64'h007ed570_01552029,
        64'hffdef4f6_00947dcf,
        64'h00910afa_010b267a,
        64'hffcc0c29_009866c4,
        64'h006d3e49_ff14359a,
        64'h00024883_00142a72,
        64'hff5ff395_0178f145,
        64'h000591d5_008f6019,
        64'hff9de675_ff37594f,
        64'h00508287_01976843,
        64'h0081fb3f_014af70e,
        64'h0077ccc7_fe35d272,
        64'h00e13755_ff95f878,
        64'h003bae91_ffebcc96,
        64'h004b64c5_0029800d,
        64'h00033964_fea7bd02,
        64'hfffbc9e3_011e9ad1,
        64'hff232456_fef9c964,
        64'h005dd0e9_fe6caadd,
        64'hff010651_ffd9dba3,
        64'h000d30b8_00ad1a28,
        64'hff5a2467_01460346,
        64'hff1123d8_fe2f6195,
        64'h00cb3556_fe87efc4,
        64'hff412a9e_ff679736,
        64'h0027afec_01432d99,
        64'hffef238c_01547737,
        64'hff97538c_0070aab3,
        64'h0083325e_002a0df1,
        64'h009bd5fc_fee878a2,
        64'hff3a9b94_ff9a85d0,
        64'hff92d0aa_00a45677,
        64'hff9b9c4d_ffbbb383,
        64'h003f3e8e_fe048d13,
        64'h00fe184a_0166c870,
        64'h0001a95d_ffa83076,
        64'hffc6c4b0_ffc24478,
        64'hff70089f_0086a7ff,
        64'h006ae183_fec473b4,
        64'h0049159f_00ecaf99,
        64'hffd26000_ffe04e3c,
        64'h0080e453_00925ef6,
        64'hff2816ff_0134ea39,
        64'h004e2c22_01bf2f7f,
        64'h009045c3_002bae3d,
        64'hffa10c84_017ba6b2,
        64'h003e3cb9_004cdf2f,
        64'h004e64a7_00ca3b87,
        64'hff22d103_0086c50d,
        64'hff3f01e7_0127a733,
        64'h00dd747a_00b02414,
        64'h002b5af4_ffb6cd45,
        64'h00a0d15d_0096c656,
        64'h00314938_014dd495,
        64'h00ed555b_fe37b472,
        64'hffd33b78_ff77f93f,
        64'hfff9cd62_fe873c6b,
        64'hff602eff_01f07918,
        64'h0017b335_fe4da8fd,
        64'h00c5dc69_00856730,
        64'h00fc36d8_014e869a,
        64'h000b979d_00c850a2,
        64'hff7219a0_fe799f00,
        64'hff290b1f_fed58195,
        64'h0016ccb1_feb1cb16,
        64'h00f20302_fea53def,
        64'h002968d7_01c197ee,
        64'hffa9c18f_ff82c9a8,
        64'h00efac8b_fe1062d9,
        64'hff7f63d4_fe9d12d4,
        64'hffc954ed_fe5721f3,
        64'h00edd12d_015cd4a0,
        64'h00ef01fb_fffa2d24,
        64'h00fd3f27_fee61eaa,
        64'hff19604b_008276c2,
        64'h002138c9_fff37926,
        64'h00ee7334_ff60c06d,
        64'h00397dc8_00f36efd,
        64'h00fcc917_ffb2d81d,
        64'hffacaa43_fef1a603,
        64'hff3dbb79_00e2206a,
        64'hffee9a81_0120054a,
        64'hfffaec2f_ff733bce,
        64'h00353d2e_fea55ede,
        64'hff355f8d_0043bc76,
        64'h00244afc_ff9ce9b8,
        64'h00516b3a_feda077c,
        64'h00c4b319_fe1c453c,
        64'h0033f867_0195782f,
        64'hfff78ba5_0161a9f7,
        64'h00b9da96_01b5e716,
        64'hfff4a7ab_00d01fc5,
        64'h00620bd6_ff853eb9,
        64'h00df85ae_01ce0840,
        64'h0001ad48_0076b400,
        64'hff065935_ffad4bf8,
        64'h004efa06_feaa1473,
        64'hff5ce160_fe10e2b6,
        64'hff9ae38c_01489d68,
        64'h00e70032_01c13699,
        64'hffb37606_fed5d74a,
        64'hffb5d1e1_ff3bbf24,
        64'hffe7895e_ff2f9750,
        64'h00bbaccb_019c495a,
        64'hffe33c97_0138258d,
        64'hffc99087_feb3537b,
        64'hffc8df93_fef32034,
        64'hff668184_003b35b8,
        64'hffeef209_002c4563,
        64'h001784a6_fe846272,
        64'hff28ba7c_ffe48681,
        64'h00289308_00cbc66d,
        64'h006c5b1a_fe100905,
        64'hff0771f0_fe0cb939,
        64'h000ca0e9_ffe67ad8,
        64'hff1e622b_011db07d,
        64'hffb49923_ff96fedf,
        64'h009a2e15_005beb26,
        64'hffa63797_008790d6,
        64'hffc8a5f8_fe7d518d,
        64'h0044cb94_ff818613,
        64'h00694e50_00d819e7,
        64'h00cc24ba_ff7f75c9,
        64'hff09bd7b_fe88bb39,
        64'h0002e9ce_01e2ae39,
        64'h00bcd900_fff22e03,
        64'h00fb25a2_011d2307,
        64'h008860a1_001dc49b,
        64'hff820ca4_fe9505aa,
        64'hff7f7d23_0058171d,
        64'hff793adf_01e853ba,
        64'hff76109a_feae9c53,
        64'h00b9799b_00f2b69c,
        64'h00dfd015_ff07a6a6,
        64'h007c92b2_0055a154,
        64'h00b61e58_00395e99,
        64'hff2f9dc5_ff581609,
        64'h00527a8c_01eea3b4,
        64'hff6dee7d_003b29c9,
        64'hffc8853e_fe3cc65c,
        64'h00d4e45c_01db961e,
        64'h00a60023_fff4ff94,
        64'h00ceba91_fe0d24fe,
        64'h00abc602_ff3f3e7d,
        64'h0082e1e3_01577b75,
        64'h0031c04c_015fe58a,
        64'h00c3ef15_004bafe3,
        64'h0029229a_ffe4c7ab,
        64'h0051d266_ff18289c,
        64'h005f4b47_019ef0d5,
        64'hffb5222f_ffb5ce39,
        64'h00ff51b7_ff41f2bc,
        64'hff6b6ce3_ffecaea7,
        64'h00506f97_fe45f06e,
        64'h0042e273_fe604289,
        64'h0076e4b2_ff4d5524,
        64'hff285c40_012a05b2,
        64'h00a5849b_ff9ed22a,
        64'h00bf3428_ffea7d7c,
        64'hff115213_fe4972ef,
        64'h00f574c4_ff35969b,
        64'h008d0498_017d5071,
        64'h0088c2bf_01ed8898,
        64'hffac9065_00ae4e67,
        64'h00d14665_01f2944f,
        64'hffd02dec_00cd9cfa,
        64'hffb6168a_ff9815df,
        64'hff57e095_ff8112c6,
        64'hff36476e_ff3bb638,
        64'hff3cbeb4_00116b90,
        64'h001a3c46_019f11fc,
        64'hff598295_01030217,
        64'hffb188b3_ff9acc15,
        64'hff306675_ff0734fd,
        64'h0023f0e9_00c677d6,
        64'hffe687aa_ffd28176,
        64'hffe94dc4_00b77f28,
        64'hffa5952c_00901696,
        64'hffdb3417_ff9c619b,
        64'h007da8f9_014f2690,
        64'h00d6c427_fea7ff6f,
        64'h00d7879c_fe63ef31,
        64'hff5567a2_00147b72,
        64'h0038a252_01770eb8,
        64'h0045dbf2_fee2dfe6,
        64'h00bc9daf_fe42e0ac,
        64'h00808884_ff380842,
        64'h00e76c2d_00ea79b9,
        64'hff647ba2_fe81d6cc,
        64'hffe4e2ee_ffe22552,
        64'h008d4369_01a18191,
        64'hfffc0684_01747675,
        64'h000073b3_011d6c87,
        64'h00e74a1e_fef62713,
        64'h00d2ccce_ff0cb7ed,
        64'h005ede26_ff373f18,
        64'hff364eef_ffa59ffc,
        64'h00a74407_fec59858,
        64'hff89997e_00ce8fee,
        64'hff059e94_fe6bc593,
        64'h00489997_00178734,
        64'h00a7fb97_00bb689c,
        64'hffe5ac2b_018773c8,
        64'hff05d0fd_febc8c27,
        64'h00884414_feb3f338,
        64'hff7b1a90_0098a932,
        64'hff5543c0_ffba0646,
        64'hff5edfc8_01a1df77,
        64'h00b523ff_ff5720ad,
        64'h00d9b510_0191cfd4,
        64'hff9bc895_0078df8e,
        64'h0068d792_ff270ead,
        64'hffb85392_fff731be,
        64'hffa6f557_01b1beee,
        64'h003a6e73_ffb144ef,
        64'h001d8d23_fe0bf9ae,
        64'h00229347_ffa13a2d,
        64'hffbb1215_017f8188,
        64'hffc250e7_ff805a35,
        64'h00b8324b_fffbdc41,
        64'hff7d2c3c_01830ffa,
        64'h00bca59d_ffdc0198,
        64'h0074f12d_010fb875,
        64'h002c3e39_00616ced,
        64'hffc8296f_00050956,
        64'hffca241f_feda9156,
        64'h004e60d7_fe11281c,
        64'hff33a5ff_ff7c93a3,
        64'h003db65f_00bec126,
        64'hffc07c97_ffb0caec,
        64'h0031f07c_011b119e,
        64'h003328a0_ff4b80d8,
        64'h009a5aac_012e6644,
        64'h00009142_01c6a89b,
        64'hff5dd8a7_004a7f42,
        64'hffc6de09_00ad85df,
        64'h00015982_01500dbe,
        64'h00f9bbf4_fed4bd22,
        64'hffb3eae3_01e73e7b,
        64'hffabe4dd_fe4185b5,
        64'hff0e06c8_01e82b6b,
        64'hff0b3aba_fec53395,
        64'hffc23161_0127896b,
        64'h00992fdc_010ece09,
        64'hff63ca6b_fffe79f3,
        64'hff951116_fec61c47,
        64'hff595810_fee419bc,
        64'hffbddd71_ffff0353,
        64'hff31a238_feac22dd,
        64'hffb339f2_feffb44c,
        64'hffac7275_fedb6b22,
        64'h007f9962_00cf9b71,
        64'h00611eee_00ea8a37,
        64'h00cd57a5_001946b1,
        64'hff76990a_ffe63247,
        64'h006a5a95_003362b3,
        64'hff7a772c_008444d5,
        64'hff8a1ae8_01850973,
        64'h00b631be_006307e1,
        64'hff11a379_fed7c2dd,
        64'h00d27b42_fff0fffd,
        64'hff79c60a_00f06ead,
        64'hfffc5a47_ffa16f13,
        64'h0005349b_fedc9d11,
        64'h004c13a8_fe71627d,
        64'h00aa2018_01f298a3,
        64'hff74729a_ffdfa8e1,
        64'h00a475ed_00170be7,
        64'h009d58bb_ff3dbe47,
        64'h00ad5128_fe58eb3c,
        64'hff754564_ff2c1d84,
        64'h0010c5db_00a6dd10,
        64'hff40a45f_01108b07,
        64'h00c12feb_00ad8ea2,
        64'hffb6abdd_fe3399ba,
        64'hffbaa42a_fe47e7d1,
        64'h00989fb8_004c3c76,
        64'hffbb600e_01a2736c,
        64'hffa3cfc7_01a22eda,
        64'h00dd9da9_fea4d9d9,
        64'h00e611ee_fec3c7e2,
        64'hfff41c23_fee76fe0,
        64'h00352891_005eaa51,
        64'h0064d0d2_0134d643,
        64'hfffb211c_ff3658cf,
        64'hff89b4de_fe3988d6,
        64'hffb594dd_0103a3fe,
        64'hff3b647b_00326cc9,
        64'hffad7d1e_ffe285e9,
        64'hff5880c4_00cbbd8f,
        64'hff9cef7e_00ad1f13,
        64'h00783307_0008edae,
        64'hff65d3f6_ffb1347a,
        64'h00283c46_fe95903c,
        64'h009264a8_ffccc87a,
        64'hffce90aa_0181345f,
        64'h00b6d187_000b7fbe,
        64'hff67b361_fff79571,
        64'h0055dc2e_fe35dcf2,
        64'hff86e845_ff1a406a,
        64'h00e403a6_fe511579,
        64'h00f66e3b_fe3df8d6,
        64'h00c2ffb3_ff3d90b8,
        64'h00a63516_01393059,
        64'h00eb7623_fe5c7cd6,
        64'h008c0afd_ffe64df9,
        64'hff957562_fe6e075c,
        64'h00105e44_0056971d,
        64'hffa93500_00a2509b,
        64'hfff04d96_ff4fb813,
        64'h009ff66a_fe38966e,
        64'h00c2e488_00113372,
        64'hffab01d8_fe22a9ad,
        64'hff674cae_019dc880,
        64'h007b26a2_ff2458c4,
        64'hff31f08b_fef65d0f,
        64'h00ef35f5_01a1c4c5,
        64'h00cf9c95_00204af3,
        64'h00b94f46_00b175b4,
        64'hffd04698_0054f8a4,
        64'h0067f52e_fe32d3c6,
        64'h008eed7c_ffdda82b,
        64'hff94093a_ffd2e769,
        64'h0033c85f_fe78821f,
        64'h0081e1a1_00c4833c,
        64'h00d686ac_ff779256,
        64'h0047eb0b_ff98ef5f,
        64'h00c5930c_01be105a,
        64'h00b69d52_fe79c418,
        64'hffb19a2d_00d44e4d,
        64'h007202a5_feb9c868,
        64'hffe12fb4_01930b77,
        64'h0077781b_ff11e47b,
        64'h0054ceab_013902dc,
        64'hff1ce0a7_fe74f75d,
        64'h00a6f6a3_fe67e6af,
        64'hff89d666_ff219115,
        64'hff025b43_ffa4704a,
        64'hff775d9a_00deeae3,
        64'h0002e26e_0057646a,
        64'hff3b9eec_01608d24,
        64'hffc3c66c_ffe016c6,
        64'hffee4c63_ffadca29,
        64'hff14e5dc_01ec4f48,
        64'h0023fa81_fece8d49,
        64'hffabfca7_ffaa7522,
        64'h001ae8e0_018bb313,
        64'hff859d15_ff361f7d,
        64'hff975432_005066b0,
        64'hff1f0e1c_01bbb175,
        64'h00b88303_fed494e5,
        64'hffb1d1d9_003cb583,
        64'hffe7a1c2_fe531491,
        64'h00167107_ff7f6c45,
        64'h003e6e05_ff2182ec,
        64'h0062414d_01e2867d,
        64'h0005e786_ff96f613,
        64'h00cf651e_fe1874e4,
        64'hff99331d_0093bbf4,
        64'hffd463ac_ff8e052b,
        64'hffb1cde1_ffbe5f9e,
        64'hffae3f2e_ffb6400e,
        64'h00ed9e75_01423460,
        64'h0076b1d7_fe8c732b,
        64'h00d56ec5_feab2617,
        64'h00de95dd_005fd682,
        64'h00c7d657_01c683cd,
        64'h00d0a407_01ff09b8,
        64'h008be063_ff465cf8,
        64'hff00ee4c_fe3019d5,
        64'hfff689fd_fe0eba11,
        64'h00b67f08_ffa95d3c,
        64'h007f5d6f_0041d5da,
        64'hff205616_019b5a7b,
        64'h00130031_014d1dfa,
        64'h006d2392_ffe7fd65,
        64'h00e6bedf_fe824101,
        64'hffffbfb0_ff06aced,
        64'hfff134a1_00764113,
        64'h003b7d25_ffc85b60,
        64'h0054dcfa_01576157,
        64'h0072fd19_00acae43,
        64'h00a40484_fe912f7b,
        64'hff4238e4_0111a1c3,
        64'hff8e6e50_ff0321c8,
        64'h00b042fb_01f6953b,
        64'h004fa12b_ff1d2313,
        64'h0001d7f2_00e70474,
        64'hffa58902_009c0a41,
        64'hfffb9260_0165acb2,
        64'h00043e4f_ffc5fe68,
        64'hff65cc9e_fff8c29d,
        64'hff650a02_01b3f812,
        64'hffde23d0_ff78d29c,
        64'hff32af1f_ffdec330,
        64'h00e54b35_005786fd,
        64'h00f2939a_013cff9c,
        64'hff18b1db_fe303a91,
        64'hffb46c73_fefde0d9,
        64'h00471793_feac5cd2,
        64'hff0d8c4a_ff2e747d,
        64'hffb99e34_ff054151,
        64'h00092e23_0108bd3a,
        64'h0087dd31_ffd2f773,
        64'h003d94c8_00ef019c,
        64'hffb20915_004feb9b,
        64'h00ca7169_0066caf1,
        64'hffe4c212_01f1dbb9,
        64'hff36f505_00bb4a19,
        64'hff94e682_00915484,
        64'h00eb3183_fe7b1327,
        64'h008a6c77_00fbe5d9,
        64'hff3c7031_006107e8,
        64'hff81a9bc_01d7de81,
        64'hff85514e_ff9465a6,
        64'h00f108b6_01f83eb1,
        64'h00c6381c_fe5d400d,
        64'hff1f1a47_fe15aca0,
        64'hff2ceb8d_00dcb9e1,
        64'h00971098_fe5d6263,
        64'h00d20cc0_fe1f55d1,
        64'hff9b91ee_ff956c2d,
        64'hff913c8d_ff9c3938,
        64'hff5e3d96_ff0eac28,
        64'h00e279d0_00c9a9ce,
        64'h003ac996_ff3b10b0,
        64'hff841a7d_fe156b8e,
        64'hff6de712_fe214850,
        64'hff9c1e51_009bac41,
        64'hffcff374_014b71c0,
        64'h003cda43_0104eb8e,
        64'h00ea3cf4_009ba9c9,
        64'h00b497ac_0153d4e4,
        64'hfff396b9_fe242597,
        64'h00c10b3c_fe561596,
        64'hffe6e91d_01a04df9,
        64'h006b4fa7_ff9159c6,
        64'h007e5761_0062e61c,
        64'h00985bb1_009d0b6f,
        64'hff3d2f39_00dce6bd,
        64'hff8a2ee6_01a45b1f,
        64'hff02b3f2_01ce385e,
        64'hfff4e0ac_fedb34dd,
        64'h0009d102_00a4ffe9,
        64'h0046d431_00cddd32,
        64'hff0919c0_fe784280,
        64'h00e01112_00f7d97d,
        64'hffa35ae1_ff71fe95,
        64'hffc60098_ffb15f95,
        64'hff2a58c5_00223e0f,
        64'hffc67bb1_fe42b243,
        64'h00899ef3_fe4f6a0a,
        64'hff838c0a_00fe4498,
        64'h00eca46c_ff372a5e,
        64'hff29e93d_fe618992,
        64'hff5ae397_ff040b9a,
        64'hff34a292_00a5537b,
        64'hffb46d2f_ffa5abd0,
        64'hff7045b7_01bdb5e8,
        64'h00366950_fefbc177,
        64'hff3fbc63_ffcb0bfe,
        64'h0039e62b_015f8463,
        64'h00a710d2_ffcdd9c0,
        64'hffc82ae1_ff62fa4a,
        64'h00135954_ff321db9,
        64'hff138bb3_ff3863f6,
        64'hffb91522_fed84d6d,
        64'h00d13b70_00d0a06b,
        64'h0030d381_00f410ce,
        64'h0021083b_01d5fcdf,
        64'h001ca2db_fffe6e92,
        64'hff5b01d2_fe3efcb4,
        64'hff8116cc_fe67451b,
        64'h0005ca50_00de6caa,
        64'h00f72d98_fea53031,
        64'hff59bd19_ff8a1533,
        64'hffb52563_ffd7e5be,
        64'hffb0e6b0_004d87df,
        64'h008d9fcb_00b61575,
        64'h0090717e_011de018,
        64'h00cd0f31_ff7516c4,
        64'h00a4c936_ff239bef,
        64'hff447c83_fe1a2326,
        64'hffaa5543_ffb8245a,
        64'h0095c3ec_017c2791,
        64'h00c3eca8_fe1e18c8,
        64'hff6d5c31_01d62455,
        64'h00d5eb29_01c61903,
        64'hff0ecf4c_00ebb079,
        64'hff6fa331_017092a7,
        64'h0029289c_fe2e2182,
        64'h00d2f2de_00b20477,
        64'h006ec37a_ff784a3e,
        64'h003f4c5a_00f1ed7a,
        64'h00813ca9_fe0fb073,
        64'hffbeb6ff_0001266f,
        64'h0020f258_ffa4af9a,
        64'h00ea663b_fed0352c,
        64'hff6697f6_fe7ff163,
        64'h00412ef6_fe81404a,
        64'hff4f6349_ff4c5db0,
        64'hff6c025d_feb79e5e,
        64'hffacf9ab_0165c1fe,
        64'h00bcbe76_0156e148,
        64'h00a73747_fedc088a,
        64'h00d21e35_0005eae5,
        64'h000ace1e_fe630701,
        64'h00ba2116_01427b50,
        64'hff0ac95a_ff68d593,
        64'h00c1071b_ffb04ed3,
        64'hff7364bb_feb5ae90,
        64'h001634c3_ffa0acfc,
        64'hffefbabb_ffb9dada,
        64'hfff47bd8_ffddc09c,
        64'hff2ace29_011052cc,
        64'hffdf478b_ffb2c564,
        64'h0088f7f0_00e19a77,
        64'hff2d6698_013cbb36,
        64'hff42abcd_ff3353e3,
        64'h0041a80f_01c25a96,
        64'h00d7df53_0044a603,
        64'h00bd035e_fe9d8081,
        64'hff2f9f3c_ff1ea732,
        64'hff820306_ff89db9d,
        64'h00a7536e_00ca0a0d,
        64'hff6d3584_ff93749c,
        64'h00781277_ffcd74a9,
        64'hffda1931_fe1c3cbb,
        64'h00d1fa05_ffb69540,
        64'hff7fd062_ff26271b,
        64'h00f42bd0_01528a1a,
        64'h00e62a0e_fe695dff,
        64'hffe8a02f_ffc103de,
        64'h00e2af09_ff4f3072,
        64'hffe02e33_003fa2a4,
        64'h0094f2cf_fe0824e9,
        64'h001a1c88_01512b3c,
        64'h00568d66_01eb26c6,
        64'h0084dc09_ffcae01e,
        64'hff5d89df_00dee01a,
        64'h007d43ef_fe4735c8,
        64'hff4a5240_013f9c37,
        64'h00422530_ff5fcd10,
        64'h00683743_01c512f7,
        64'h0016ffc1_fe328a11,
        64'h0071305e_fe09404f,
        64'hff833e89_01e4fbd0,
        64'hffa320d9_ffe677b8,
        64'h001bb72a_fef925e9,
        64'h008931f2_fe79a1d5,
        64'h00629793_0069f1dd,
        64'h008598ef_00327cf1,
        64'h004bf927_ff6cde4f,
        64'hff1740cb_fefffe19,
        64'hff426907_00325951,
        64'hff5ecab1_fe8efefa,
        64'hff5973ce_fff24859,
        64'h00c1a16d_ffc76bad,
        64'hffa78a6b_ff1dd3ab,
        64'h00c63236_01393a9b,
        64'hff0f7a3c_01b6368c,
        64'hff996f80_00e274c6,
        64'h001ef4a5_00a200f2,
        64'hffcbcc76_00394627,
        64'h00399164_012219f7,
        64'h0065cdce_00a2a1a5,
        64'hff220c8c_fef27dab,
        64'h00238e6c_ff82b1f5,
        64'hff1ffe0d_ff62127d,
        64'h00e8e914_00f63a30,
        64'h00b9be7c_01c5f0d0,
        64'hffe7977c_01f533a8,
        64'h008f570e_007c1853,
        64'hfff98002_00bac89a,
        64'h00775591_004725fd,
        64'h00b5cc96_001d6193,
        64'hffb73b96_00c8d4f8,
        64'h00af808d_017b2c0e,
        64'hff4de0dc_fedfe111,
        64'hff9be032_013a637b,
        64'h00c0e33f_001b3276,
        64'h00b5b9b7_fff04f06,
        64'h003e3f8a_ffec2847,
        64'h00975197_feb3e1cc,
        64'hff42f722_ffdc8e5c,
        64'hff04fa96_017441dc,
        64'h00e55366_ff7baf14,
        64'hff62b8d2_0108589c,
        64'hff3eda97_018bd093,
        64'h004f120e_fe799c59,
        64'hff4b930e_01d72b21,
        64'hff347651_00c0955f,
        64'hffdd3be2_fee35288,
        64'hff9ad417_009dc9ec,
        64'hff9a6996_fe457089,
        64'h003a9c48_0017d489,
        64'h00c55fa8_fe2e7422,
        64'hff6a84a4_00338b0f,
        64'h00440419_01c23d6b,
        64'h00695bef_fea62ba0,
        64'h002677b0_018e71a5,
        64'hff13ee21_ff5ceae7,
        64'h00ef3cce_0186c60f,
        64'hffad78df_01f58c52,
        64'hff573c7b_ff62d550,
        64'h0062eb7e_fe70a5b8,
        64'hff18683f_0127923d,
        64'h00794990_015b12fd,
        64'h0031c4a8_fe062b62,
        64'hff82d8f0_febf508a,
        64'h00e5bf60_016997e6,
        64'h00baac5c_018830d4,
        64'h0002f2c6_0020568f,
        64'h002f4789_009dd1aa,
        64'h00c7a0ed_00161d08,
        64'h00383a76_006d24d3,
        64'h006bde53_01a86c34,
        64'hff4cb235_0191669e,
        64'hffaedbf0_01cc5ad0,
        64'h005081a1_ffdb54e5,
        64'hff9a5c0a_ff661df0,
        64'hff273b5e_00f297ef,
        64'h00ca0aee_00f713ad,
        64'hffcffec5_ff986864,
        64'hffcda79b_fe92493a,
        64'h0037f3bf_fea53320,
        64'h005070b8_011f2622,
        64'h00e64285_feccf20c,
        64'h00acb836_011a78cf,
        64'h0096c9a6_ffbd2680,
        64'hff3c8e00_00cabb77,
        64'hff86a0e7_011fb576,
        64'h00b1e428_ff667c20,
        64'h00510d37_00c5caed,
        64'hffa68664_fe64f1ce,
        64'h00e2c141_fff3d8f1,
        64'hff834030_0170ecb7,
        64'h00b5fe53_00e94386,
        64'hff114978_ff200d6a,
        64'h00a4e1ef_00d14eb6,
        64'hffe80e56_00d3f966,
        64'hffe5cadc_00397b68,
        64'h0008b482_fe60684d,
        64'hff497b68_fec4e5f9,
        64'h004196ac_fe50d8cc,
        64'h00b76491_0061c62b,
        64'h0029ceba_01f079fc,
        64'hffc1c95a_010a8428,
        64'hff1ba9fc_01498140,
        64'hff1b3d31_0073daf0,
        64'h0039e897_01714088,
        64'hfff6c483_ffcf92ab,
        64'h009c36ed_019afb76,
        64'h0057614b_fe18188d,
        64'hff87f3bd_fe658fc6,
        64'hff3242bd_01c7f107,
        64'hff7f7b0e_01f1b278,
        64'h00315aa9_fe2c1c92,
        64'h00bcb82d_ffb2a237,
        64'hffa1a609_005d352e,
        64'h0007b655_01544690,
        64'hffb6a631_ff8d5572,
        64'h00fea4a0_013a8be6,
        64'hff888602_fff8f59f,
        64'hffec77d3_ff73890f,
        64'h0086d051_008e333d,
        64'h0094f0f5_fea50881,
        64'h00239467_007e2b3e,
        64'hffb37e4e_010be1e3,
        64'h00b2d9c6_ff4ff60a,
        64'h002fde46_ff6fd18b,
        64'hfff5585a_00df4f5d,
        64'hffd33ad3_ff7d1175,
        64'hffbaf348_ff0db188,
        64'h0088540e_fe03d8c2,
        64'h00b32f3f_012c9235,
        64'hffd7036d_ff7528f9,
        64'h00bb5336_015659a6,
        64'hff09c2b1_003d6954,
        64'h009e9b20_009ae5d3,
        64'h00821894_fe7a49b6,
        64'h0082438a_ffab3119,
        64'h0030c367_00a11694,
        64'h005572ca_00d18df2,
        64'h00c98157_00f5b277,
        64'hff785606_fe177130,
        64'h003dea34_fe827b42,
        64'hffee0bd2_feb3bcab,
        64'h00c78662_00bb79bb,
        64'h000ad358_fe242941,
        64'hff2c8052_fe886eeb,
        64'hff4f9568_fe53f9c5,
        64'hff300060_fe8f632a,
        64'h004f62db_00951364,
        64'hff0ec987_01c9aeb5,
        64'hff0b311a_0112c10f,
        64'hff09357d_ff8117ac,
        64'hff82a564_01839e9e,
        64'hff1d9240_ffd4ce32,
        64'h007492a2_fed83741,
        64'h006313c2_ff0a290f,
        64'hff5a5572_00ce15a3,
        64'h00ab75ca_ffa806c5,
        64'h00ae78fd_013533eb,
        64'h000ea8c5_0107e1e5,
        64'h00ea8f93_01c2c8ec,
        64'hffa14f5c_0018a9af,
        64'hffbb111c_00d72262,
        64'h0034db30_019d3bb2,
        64'hff5af6bd_fe38db41,
        64'hff958cde_009dd3f4,
        64'hffc9316b_ff5a51f1,
        64'h00de51bf_fe4b5f07,
        64'hff1d2717_ffa295b3,
        64'hff0f8851_fffbc1de,
        64'hffc0e58c_01e631d7,
        64'hff86cc52_ff3cc76d,
        64'hfff63a64_01b5569a,
        64'hff87f537_01ba91af,
        64'hff8902ab_00ebaf73,
        64'hff4d82cf_ff4bd6d0,
        64'h0081f931_001a54bc,
        64'h0065e968_01873e86,
        64'h008b5992_00f940cc,
        64'h00241342_ffb8777a,
        64'hffcbd671_0023de76,
        64'hff401260_0183fa2a,
        64'h005b63ec_01534c47,
        64'h0076f01c_00cdd196,
        64'hffd6e8ee_ff97fac4,
        64'h0000fbc4_fe2d70b1,
        64'hffbbfd85_fe53c90a,
        64'hff833842_00a925f1,
        64'h00c56e41_0170a2a7,
        64'h008b5822_019a6259,
        64'hff90d4b4_feaed289,
        64'h0060cde4_ff7f146a,
        64'h00719f02_fee6210e,
        64'h0013237a_00efd13c,
        64'h00fa3fa1_ffd032f0,
        64'h0026f5f4_00feaee3,
        64'hff412644_fe410cec,
        64'h00167c6f_00877507,
        64'hffa3c08e_009e5fc8,
        64'hff8ede58_ffc7ad32,
        64'h00aba38f_ff836c8c,
        64'hffa8f909_fef22d87,
        64'hfffa7c28_fe79652e,
        64'hffea7167_002ec4f1,
        64'h001e8654_0152e096,
        64'hffd15a30_fe1781ac,
        64'h00fce461_fe97467d,
        64'hff860124_00cd7ab3,
        64'h0018e705_feddb0a4,
        64'hffdecb90_ff05d3ea,
        64'hff35fbe2_009b621d,
        64'h005b9840_fe7e6a4d,
        64'h00f090e7_015f3e22,
        64'hff25ace0_ffdfbb41,
        64'h004c61bd_ff1e3929,
        64'h00b91718_feb4938b,
        64'h006385dc_fe399ffe,
        64'hff5a225e_ff966aea,
        64'h000ad2cf_ff144951,
        64'h004ba640_0086e4fd,
        64'h0087a969_00fca45f,
        64'h0030f7a8_fe314e89,
        64'h007c903d_fe253126,
        64'h0051eacb_ffbea455,
        64'hff451178_014ddcd5,
        64'h005e9846_fe5eee37,
        64'hff6b2600_0105efcf,
        64'hff3ccbdc_ff723297,
        64'hff89797c_0155c1c6,
        64'hffb7b018_fe34aca0,
        64'hff6006af_00a11229,
        64'hffb8ea43_fefb8d0c,
        64'h00f3102f_00a460a1,
        64'hffbb3919_00fa7012,
        64'hff9da303_017317b9,
        64'hff598795_ff391ffa,
        64'hffc3ef49_fe6bdda2,
        64'hff6dd81b_fee779bb,
        64'hffb35430_00d5d069,
        64'h001e705c_00bd843b,
        64'h0071036a_01ed3c06,
        64'h001112fe_fff30fde,
        64'h002983e4_018d61a5,
        64'h00250994_0066e80d,
        64'h0094a97d_fee81ed9,
        64'hffee1935_ff150933,
        64'h0009167a_0165f0e8,
        64'h00a2ab38_002e9d9e,
        64'hffa8bbd7_01a27ae1,
        64'hff256019_00e83c56,
        64'hff0142dc_0095afdf,
        64'h005b8726_00746d9e,
        64'h00f7b966_00b1f200,
        64'h00d1c133_009d28da,
        64'h00560f5e_ff83c1cc,
        64'hfff0c153_ff0a1c5e,
        64'hff51e2f0_fecb4f0e,
        64'hff1ac479_01c7d818,
        64'hffc76542_0042a94b,
        64'h00001f58_0097bd3a,
        64'h00b78ca5_ff241bb3,
        64'hff581e31_fe43a923,
        64'h000e34fd_ff5b95f3,
        64'h00183321_fe59838d,
        64'hff763962_01ca1003,
        64'hffd3a4b2_011838f5,
        64'hffaaa3b4_01537ebf,
        64'hffcf0be7_0032d6f6,
        64'hff85e5ac_00dbf106,
        64'h0018878b_007d3305,
        64'hff0f8420_00a7f3ba,
        64'h004ce02a_ff2f031d,
        64'hffe15af0_fece2d26,
        64'hffbc5025_0022e51a,
        64'h0070f416_ff75d0ee,
        64'h00cdf218_01db00cc,
        64'h0082e396_00f9870f,
        64'hff09c1c1_0033701a,
        64'h0094e9af_00cba34a,
        64'h00e1d431_ffb66d13,
        64'hffcab693_feb54f0c,
        64'hffc70990_007eec8c,
        64'h00e895e7_ff0fd9b5,
        64'h001bd008_016bc059,
        64'h0070d483_fe35ea65,
        64'hff76c1ab_ff9215ee,
        64'hff1fc1c0_fe2819ad,
        64'hffd70f76_005370ff,
        64'h00fee72f_0008dd12,
        64'h001f5e72_ffe8beab,
        64'h0021b66e_fe18b637,
        64'h0042b83d_ffc8722e,
        64'h00dd8239_ff60d1a7,
        64'hff5ac8f1_ffd330b2,
        64'hff1edfff_0125dd40,
        64'h008a59cd_00cc5fb7,
        64'h000b1ec5_0160fb43,
        64'h0079edbb_00d4fafe,
        64'hffe4eec2_ffaf9766,
        64'h0003e501_011ee040,
        64'h00a86f69_016ae6e9,
        64'h004a88ed_fe936bc9,
        64'h0048a1a6_01b7aeca,
        64'h00c17681_ffdbf7e5,
        64'hff6a74ba_00c2733a,
        64'h00699fb4_fed75302,
        64'hffefde03_fec540a8,
        64'h00591a28_01dc24d3,
        64'hff482326_ff810862,
        64'h007fb9fc_0000fe06,
        64'h00870791_fef3cb94,
        64'h00d04450_01eaa936,
        64'h0032fb2b_00de00fe,
        64'h00fd8d75_ff2a7627,
        64'hffcb91ca_0130f317,
        64'hffbf5eeb_01dde6b3,
        64'h00d94b36_01706ffe,
        64'h00a12884_ffb42d5e,
        64'hffeea7cd_0052869b,
        64'hff513525_fe92fc86,
        64'h0027d5a4_000584fe,
        64'hff3a17b2_003e5255,
        64'hff81febb_008306fb,
        64'hff94fec7_fea731a9,
        64'h00a00180_fe6c8341,
        64'hff82fb94_00c4b627,
        64'hffe5bae6_fe3642e0,
        64'h00361692_00c0845a,
        64'h00abfd4c_00976b86,
        64'h007fbc94_ffa800f0,
        64'h00616236_015dc389,
        64'h0017170a_ff7498bc,
        64'hff0155a7_01cf475f,
        64'hff57037f_01f05d96,
        64'hff2c3b9b_0021c58f,
        64'h0098df9b_00bd64f7,
        64'hff847b3e_ffa7d411,
        64'h00f7fb82_ff737868,
        64'h00c6b791_013f0caf,
        64'hff854702_01fa131b,
        64'hffcae996_00bcda9a,
        64'h00eca7a0_fe6c66f0,
        64'hfff0a9d6_fe92f2f6,
        64'hff0e5d98_00e668fd,
        64'h00143b29_012651e5,
        64'hffc71fc5_01c2ecab,
        64'h007197f5_01c6f262,
        64'h00d82b33_fe580a32,
        64'hff6e59fb_fef93ac5,
        64'hff0f539c_0112cd40,
        64'hffa000b7_015eaba9,
        64'h00f733de_00c385c3,
        64'h0014ca45_ffb7ba98,
        64'h00202423_fe182fe2,
        64'h0080287a_ffe382f6,
        64'hff036714_ff1d9316,
        64'hff8906c3_ff0ebc49,
        64'hff3d299e_ff3b0ba9,
        64'hffaf1143_fea4d801,
        64'hff5d7ba5_fea4a0c0,
        64'hffeace56_016f9a4c,
        64'h00102199_01656429,
        64'h0014b686_01b850aa,
        64'hff97b997_ff167bff,
        64'h000e31e0_ff684817,
        64'h00329da8_fe789686,
        64'hff356481_fe10e591,
        64'hff19ed4b_ff561c72,
        64'h000e9477_fe300df4,
        64'h007bd3ec_01594706,
        64'h006d7aee_fed631e9,
        64'hff085475_002a822e,
        64'hffc3bfb2_ff2a5e79,
        64'h007b6029_fed54245,
        64'h001e6fea_01b08792,
        64'h008276f2_feb804e1,
        64'hff4fb467_fec12ec1,
        64'hff87f104_01a3eb86,
        64'h007792f3_002af3c6,
        64'hff23ba6e_ff8693a0,
        64'h00a57686_ffb400db,
        64'hff8cd331_fe5dbacd,
        64'h00a84726_0119f2d5,
        64'h0010f04d_01ee1fd7,
        64'h008c7e5e_01bc6f9b,
        64'h006ab219_019e371e,
        64'h00efe931_01da6dc9,
        64'h00add5e5_01ec05e3,
        64'h00123739_fe4baec6,
        64'h00d8fa66_01ddd97c,
        64'hffa31ef7_fe6f4159,
        64'h00216131_fe930566,
        64'hff6c9d44_01755dcf,
        64'h00adb9e8_0128b071,
        64'hff5f47a8_0084827b,
        64'hff2f8877_00f970b9,
        64'hff8f453b_00db4297,
        64'h00c59f3a_ff2663fe,
        64'h00e6a161_01e07080,
        64'hffb8c603_0098b648,
        64'hffb212e6_01bb55db,
        64'h002d0695_00c6670b,
        64'hffb3c07e_ff0a8d7c,
        64'hffbbaf98_0084035e,
        64'hff824f73_00bc2951,
        64'hffcc8f0c_00026189,
        64'h00c5dd87_01d621e5,
        64'hff987f6e_ffd27b99,
        64'h00f8de8d_01444496,
        64'hff91637d_001e273b,
        64'hffd600e7_0078ea1b,
        64'h00c24df7_00b0a5b0,
        64'hff5a7bb6_fe77b128,
        64'h008bdfb8_ffb8710f,
        64'hffec1278_feca062c,
        64'h00fea7d3_0105d613,
        64'hff5c0ed9_0159a83c,
        64'hff7b058e_00339aeb,
        64'h00ab66b6_01f3c19e,
        64'h0064868c_016baebd,
        64'h0000cf00_0102c086,
        64'hffadd6d9_00a66099,
        64'hff090b08_01364dca,
        64'hfff78045_01f65be5,
        64'h00fc2eb1_ff91d313,
        64'h00805775_fef6ef49,
        64'h005c77fe_fe8c575e,
        64'hff79e376_00ee29dd,
        64'hff04b2e6_000df999,
        64'hff42bdec_fed84afa,
        64'h00102332_01469954,
        64'hffc86aae_fff4e36b,
        64'h00f32240_fe02e481,
        64'h00d63371_0077a4ae,
        64'hff281f85_00e5e895,
        64'h00f98ca1_fe994ced,
        64'hff506eef_ff2cac49,
        64'h00a3963c_0006ccad,
        64'hffddfa72_ffd96574,
        64'hff6a8fb6_01d95a23,
        64'h005cd1f2_01da81d3,
        64'hff3db36e_016b8ae8,
        64'h005d6a46_0016913f,
        64'hff41628e_002b3406,
        64'h006efeca_004e98f8,
        64'hffa9da5a_ff5530b1,
        64'hffb7a023_017ab1c8,
        64'h009ae46d_01ae44f3,
        64'h002abe6d_00b75601,
        64'h0084e638_00ca1635,
        64'h007face1_01cac65a,
        64'h00bd42ed_ffcf0c15,
        64'hfff2fd6a_fe3b16c8,
        64'hff474d53_01296ec6,
        64'hff83e9fc_fe96fd79,
        64'hffe8583c_009f4136,
        64'hff6d00ea_ffcbebe8,
        64'h0081bc8d_00bebe1c,
        64'h009a2b18_01a73b1d,
        64'hffc14c13_ff8fb009,
        64'h0052a249_012cbbe0,
        64'h00c8d200_ffd1a93f,
        64'h00d03079_004232a0,
        64'hffb3afaf_014dd73e,
        64'hff5df853_fe34bee8,
        64'h0097a046_fe1c04fc,
        64'hffccebd2_01310da5,
        64'h00acdee1_ffa86189,
        64'h007261e0_fea52db7,
        64'hffd1b1b2_fed1d825,
        64'hffdfe9e4_00f9e584,
        64'hff73646e_00c7dc1d,
        64'hfff0ad20_ff4682fe,
        64'hffd038c3_008d3995,
        64'h0025eaf9_ff8cc8c8,
        64'hffe0bf16_01682ab5,
        64'h0099465d_003ebfe1,
        64'hff188520_fe7bb03e,
        64'h0019d5ac_011be821,
        64'hff55b472_00312ad7,
        64'h0037a95c_fe50e365,
        64'hff6b4685_fe2cd7fb,
        64'h00a48c19_fe7c2390,
        64'hff5aeed4_ff7a578a,
        64'hff9f52b2_00c343e9,
        64'h0076012b_fe8ce9a4,
        64'hffcd0edb_ff2d6929,
        64'h00a8af6e_00a86f50,
        64'hff23992b_ff0168ff,
        64'hff12b301_003241c5,
        64'h0042fa6b_0012a6c0,
        64'hff46903d_fea963a4,
        64'hffa6a426_ff1b0129,
        64'hff52dca4_fe217535,
        64'hfffc60b4_006e7ce3,
        64'hff534e3c_ff70cffd,
        64'hffa699fc_ff580c0e,
        64'hffd6455c_012c3a97,
        64'hff26d187_fef67bd1,
        64'h00d47849_01bc5699,
        64'hffc17d3e_ffb1e523,
        64'hff3d555a_ff694a7d,
        64'h0064209b_ff31f68a,
        64'hff459a4a_01dacfaa,
        64'h00bd8df6_ff491e6e,
        64'h00084fb8_010dfcea,
        64'h00f18021_01d700b3,
        64'hff3b2ae2_feac6f47,
        64'h0015858e_fe9b4dcd,
        64'h00458248_00961548,
        64'h000b2627_008b6bd5,
        64'hffb0d254_ffee2f4e,
        64'hfff7b5aa_016a6d09,
        64'h00f576a3_fff1b645,
        64'hff0e8e13_01c9e05c,
        64'hffb627db_ff2f88f6,
        64'h00224c1b_008f3547,
        64'hff15e54d_006fe8b7,
        64'hffa39f92_01c02a2a,
        64'h000b1453_ffb2a277,
        64'h00f836aa_009443bb,
        64'hff0d35cf_ff60c8a1,
        64'h004c9ef4_001c2668,
        64'hff2d44d5_feb434f2,
        64'hffd95e69_fe9e822d,
        64'h0002ddfb_fe5f78aa,
        64'h00d56feb_fe71dd17,
        64'hffe68803_ff854230,
        64'hfff6cb47_fe5d9aaf,
        64'hff18e570_ffdcadd9,
        64'h00c66ae9_018235b3,
        64'h008fd2df_ff32eb43,
        64'h005ad933_ffdd1184,
        64'hffd001c3_fea743e9,
        64'h00e549d4_016e7f8f,
        64'hffd30087_fe1fec1f,
        64'hff5d6968_fed71bdd,
        64'hff471a83_ff316c58,
        64'hff2786cb_fe416fd1,
        64'h00101297_00a0afbb,
        64'hfff874a2_fe1d3c8e,
        64'h00bc5fa4_004aed8a,
        64'h00561ad1_009e1a1e,
        64'hff054935_ff96463d,
        64'hfff1562f_011c6f65,
        64'hff0efa2b_0181397e,
        64'hffb2d290_fec89a79,
        64'hfff6dc3e_000b3a4a,
        64'hff71f41c_ff1f045a,
        64'hff69aa6d_ff0a314e,
        64'hff9078c7_01e9096b,
        64'hff5cc5ab_0035b642,
        64'hffedf0e4_01a45db9,
        64'hff20521a_01bd6958,
        64'h0030a871_00bcda29,
        64'hffb93644_ff78c5a7,
        64'h005a1365_fea0410c,
        64'hff452244_017898c6,
        64'h005ef4c8_00324ce4,
        64'hff60bd12_fe752da6,
        64'h007ee7de_0036fe39,
        64'hff3eaf1c_011055f9,
        64'hff2fa861_01efd999,
        64'hff2df1ee_fe6e1f8d,
        64'h005c0e10_018eaf67,
        64'hffeb84e9_ffd7fa3c,
        64'h00121965_00c3d89a,
        64'h00932632_febf72d0,
        64'hff153a47_00529ccb,
        64'hff2c510d_ff62d079,
        64'h00c1a084_00165c51,
        64'h009aba2d_fea9bc29,
        64'hff2cee72_00d261bd,
        64'h00af7d26_ff4c23d4,
        64'h00b9dcd9_014707fa,
        64'h00f6d612_01ff737b,
        64'hffa64807_ffeae2e0,
        64'hff77a554_003b22af,
        64'h008c5911_ff373409,
        64'h00150d86_00a01600,
        64'h004a6314_013ae9dd,
        64'h00e21d6d_fe883564,
        64'h00ba80af_003eb54c,
        64'h0080b854_fe5df981,
        64'h00b61cfb_01e7af6e,
        64'hff53eb06_01c0fead,
        64'h0076847c_015d74f8,
        64'hff2582e3_fe347fef,
        64'h00513017_00e997f4,
        64'h00d74c2a_019b4d59,
        64'h0030ae18_ff39caca,
        64'h00f0a4c0_013b9ec5,
        64'hffe76760_ff5d0173,
        64'hff261e24_01610042,
        64'h001d0cf0_fe3cb394,
        64'hff7bdc24_ff3b0c89,
        64'hffea79c7_ff788dee,
        64'hff6bf37e_ffc0d058,
        64'hff4c51d2_0112100a,
        64'h004818cf_ff4947d0,
        64'hffca9d48_febd1ff9,
        64'hffa671cb_00138154,
        64'h00bea7fa_01022efe,
        64'hff4fbbb1_ffefc57a,
        64'h00bfce78_fe85485f,
        64'h00df2b9c_01c17c5e,
        64'h0026c3a9_ff2325db,
        64'h002e622a_01c93b03,
        64'hffcde4fd_fe66c55c,
        64'h0022e9a6_feb531d6,
        64'hff7b0670_004883f9,
        64'hff2d1573_0123bbbe,
        64'h0077a963_ff3185bf,
        64'h00d6ea2e_fec2c9a8,
        64'hff637b62_fe1278ec,
        64'h003eefb9_fe0aa4ed,
        64'h00b7ca05_00c8d473,
        64'hffae758f_ff560b6e,
        64'h009761c6_0132995d,
        64'h006b88f4_feb960cf,
        64'h00ba1aa2_00e38770,
        64'hff0155dc_ffa96c98,
        64'h0041323d_ffb037ea,
        64'h0096878b_ffc9c8bd,
        64'h001b8570_fe54c1dd,
        64'hff073a78_0104e1e4,
        64'h00756afb_fec76e21,
        64'hff3ccbde_fe7a0c07,
        64'hffb7d5c8_01d34e6a,
        64'hffd174c0_ffa9c0cf,
        64'h003c0f80_ff8658de,
        64'h003135b1_fe19c6dc,
        64'hff6188d9_ff701027,
        64'h002e9947_005b2b5a,
        64'hff9dac98_008b8d2d,
        64'h00645d74_009f8384,
        64'h00455010_01855661,
        64'h00e989fa_018d52ff,
        64'hff44c565_00dfd2ae,
        64'hff082fcf_fe79b424,
        64'hff8dc377_ff43d73b,
        64'hff2ae0a0_fe4539a4,
        64'h005898f0_00c9842e,
        64'h005ec344_ff5375a6,
        64'h00b50b88_0108ead4,
        64'h00e029ee_01e64fbc,
        64'h009eaefc_001fda31,
        64'h0042b96a_fe7e42b1,
        64'hffbe8c59_ff6863c2,
        64'hff0093c3_feb59d6b,
        64'h00e7d612_017018de,
        64'hff5b6df3_fe1b9f99,
        64'hffab28a4_ffb9a30c,
        64'hffa58bfb_feb1a9db,
        64'hff99e3f6_fe9108f3,
        64'h00f84779_fffb62a8,
        64'h007031b1_ff80e5ee,
        64'h0017f745_ffefc30e,
        64'hff579314_00fe12a9,
        64'h002f32ee_ff2a2a86,
        64'h00ac30e1_013756e8,
        64'h00945111_ff34afbc,
        64'h008c4cc2_01077866,
        64'hff4d8d81_0015171e,
        64'hff2bbf40_ffb71a03,
        64'h00ca035e_003d05fc,
        64'hffd15ed8_fed9d513,
        64'hffab8671_ff78bb88,
        64'h0099ec61_ff4e246a,
        64'hff3d9d7d_0130239a,
        64'hfffb2ef6_ffe33122,
        64'hff12aefa_014df54a,
        64'hff473fb0_fffaffd9,
        64'hffef0327_ff056f98,
        64'h002b5c97_01b29ecb,
        64'h00574743_017a8bd5,
        64'h007da415_00daf29e,
        64'hff40928d_01a532d4,
        64'hffb90141_015ce6a1,
        64'h00840bf7_ffa2b20d,
        64'h00ca0124_003d0eb9,
        64'hff7af1b9_014e5f6a,
        64'h004f2bb0_fea36a22,
        64'h00e3b1e3_01f6b0fe,
        64'hff9521e3_00ba97cd,
        64'hff3f7637_ff9dde6d,
        64'h00bc06e5_01522646,
        64'h003c7d53_001e39a5,
        64'h009979de_ffd1f528,
        64'h004d1843_fe6ab7da,
        64'h00ec055d_018e9533,
        64'h006eec17_002ca1e2,
        64'h00e3372a_01b5fbf9,
        64'h0011a346_01267cb8,
        64'h00b4977c_feb256b1,
        64'h00e74483_00d7de03,
        64'h00c28bdd_00b11f8c,
        64'h00c38781_ff51cb7e,
        64'h00574a39_012bc66a,
        64'h00152a93_ff316b39,
        64'hffbba220_0078ac24,
        64'h00017973_01c7ddf8,
        64'h00a8d74f_00fcd454,
        64'hffe03c5a_000c3a94,
        64'hffe3683f_0061073f,
        64'h007d70ef_01fb69dd,
        64'hffa4de27_0186b8b4,
        64'hff51d489_fea26910,
        64'hffb65306_012fe6ad,
        64'h0048f83c_ff6b9302,
        64'h006127da_ff503c8b,
        64'h00b39637_018d18a9,
        64'hffb52191_008b4e5c,
        64'hffdcabcb_019b1d3d,
        64'h00593b4d_00b18161,
        64'h00e002dc_01273152,
        64'hff42f505_fe53867b,
        64'hff6afc88_ffd7592b,
        64'h0071b15e_0087b6ad,
        64'h005ab35e_01718532,
        64'hffaec801_fe0cbdd4,
        64'hff9ac193_00c2e08b,
        64'hff0ac913_00af353b,
        64'h00a2a84d_fe621edf,
        64'h003fb8fa_0071e188,
        64'h000111d8_fea1a1bb,
        64'h00cfbcd2_00f2d250,
        64'h00c230da_01291635,
        64'h003b45cd_fede67c3,
        64'h003474ac_ff9ffeb6,
        64'hffa2d129_feefccd2,
        64'hffba1bad_01a1ca13,
        64'h001827d3_00f2883f,
        64'h00030abd_01f85c6b,
        64'h0092ec8c_012a9952,
        64'h00913378_00dbf096,
        64'hff389124_ff0480a6,
        64'h003cc19b_fe05b5f0,
        64'h009b108c_fe3622f4,
        64'hffc00d13_fe30cd9a,
        64'hffaedc27_01f019d5,
        64'hff06d903_fe5fee2b,
        64'h001a3e9d_ff8e118e,
        64'h002539f6_ffdced3d,
        64'h00c7ea16_fe62241c,
        64'h0050c4f1_018a0fda,
        64'hffd38e20_fedfbdfb,
        64'hffb2acef_fedb9c96,
        64'hff8cee4a_006bcd34,
        64'hff05e485_01c735a5,
        64'hffe83f14_ffea6cd0,
        64'h00e4db2e_01ab20ea,
        64'hff3843c4_00da0f3d,
        64'hfffdefb9_0048cd77,
        64'h00b83eb2_fe363948,
        64'h0092b2e6_01e0f9b4,
        64'hffe09b5d_ffb8b9fb,
        64'hff4a3633_fe31acac,
        64'h00651428_ff6fec0e,
        64'h00cae185_ff816a54,
        64'hff9cbc81_00c17007,
        64'hff852564_01d094bc,
        64'h0056bbb4_002f523b,
        64'hff259f6e_00ed7e13,
        64'hffc30b76_00a7ad16,
        64'h00dcf9f5_0031186a,
        64'h003c4957_ffc2d13a,
        64'hfff3bda3_0014a053,
        64'hff00b4dc_feb419bc,
        64'h00363307_0048bc17,
        64'hfff093ff_00f8fedf,
        64'h0069b890_00d5bdd6,
        64'h0084f732_fead36ac,
        64'hffe80f8b_fed10853,
        64'h009d8dd4_01737c53,
        64'hff4aca12_ff2dce08,
        64'hffa1020f_017769f5,
        64'h00f60b2e_ff7b07b9,
        64'hffc40626_fff1acb7,
        64'hff8dd56f_013a976f,
        64'h00826f29_fe89f238,
        64'h008e85d2_fe61a67c,
        64'hffa768bc_003c1551,
        64'h00ba12d0_fec2a06e,
        64'h0042f271_ff12ccfd,
        64'hff5561ca_fe0b586b,
        64'hff3028f6_fec1ae49,
        64'hffbe4f9b_fea3416c,
        64'hff626f0f_fffd8bf1,
        64'hffc35dc9_008d9b66,
        64'h00edbdf8_fe202b5d,
        64'h00492eb2_01131da6,
        64'h00daa524_01956e05,
        64'h00f1709f_00ae6d24,
        64'hff8314bc_fef2bb9a,
        64'h009c87d6_fe5de6a4,
        64'h004f9068_ffeb1b46,
        64'h0074ced8_fe8ce344,
        64'hff21eac2_ff4eb7a1,
        64'hff1e2751_006fc917,
        64'h00465260_0067e91e,
        64'hff50f22d_0126f9f7,
        64'h00386b8e_01a9e9cb,
        64'h004853f8_0194962d,
        64'h00ad1301_003677db,
        64'hff46bb81_01ffd591,
        64'hff687892_fee37b76,
        64'hff8343f0_fe5ce50f,
        64'h00614b57_017cb208,
        64'hff7f858a_0048ce22,
        64'hfffa73fc_ffcf7290,
        64'hff8c78dc_015c9a59,
        64'hff1a5817_ff994372,
        64'h0076d264_01b42bc6,
        64'hffe56b20_00d1bf65,
        64'hff885e84_00e1c198,
        64'hffe33849_fe0a7534,
        64'hff02a633_0075a1cf,
        64'h0093ef4c_005fa0ce,
        64'hffc1166b_01b7daf6,
        64'h00eb9d64_febce4bc,
        64'h001cc7e5_01cf7f27,
        64'hffa61e0e_01ec366e,
        64'hff9c1bbf_007c3497,
        64'h00713dd0_ff2c6a58,
        64'hffe15b98_0173bea5,
        64'hff35d66a_007772f0,
        64'hff9bdab5_0003619f,
        64'h005a2166_fefc9058,
        64'hff9db75c_ffccad85,
        64'hff5ee636_ffe38469,
        64'h001e17cf_fea11c95,
        64'h005971c5_01940dd9,
        64'h00a39997_00a59cda,
        64'hff6320e0_ffa0e8a8,
        64'hff3539bf_fedc479a,
        64'h006277ad_fe6507e8,
        64'hff1f7a0c_0040c29f,
        64'hff875772_004c97a6,
        64'hff236a96_016fb925,
        64'hff555f9c_006ea621,
        64'hff0f030f_ffedcf84,
        64'hff4dd050_0065a464,
        64'h008813cf_fe156354,
        64'h00887f52_0073cf08,
        64'h006b49eb_feff1bd2,
        64'h00875151_fffdeee1,
        64'h006113af_00233526,
        64'hffcc6426_ff564ca8,
        64'hffb1452a_fe334424,
        64'h007d3a94_00fc49aa,
        64'hffddbd59_fe9afc53,
        64'h00b0bb85_009e34c2,
        64'hff6df62d_fe8a47e4,
        64'h00c5c6ca_feaaf1ee,
        64'hff9241af_01a4245e,
        64'hff477ca0_01c8ad69,
        64'hffebf872_008276ba,
        64'h00f0f462_ff978af8,
        64'hffa81c74_fe17b807,
        64'hff8061a2_01d37308,
        64'h00211e3e_fe823b62,
        64'h000653e3_ff06095f,
        64'hffd98e18_fead2d27,
        64'h004e1f11_001fd404,
        64'h004d8457_01ff295f,
        64'h00927ad4_fec18f7a,
        64'h00f623ed_008bf3ab,
        64'h009c4051_ff307a7f,
        64'h0008860d_0110be8e,
        64'hff974551_ffec52e2,
        64'hffbb588a_003cd92e,
        64'h00ecffc1_01811f2a,
        64'hff37ec69_ff05bdd1,
        64'hffd7dda4_014a3189,
        64'h00dd5ae4_fe889bc8,
        64'hff71acc1_00905aed,
        64'hffc7c4a0_fe13ad49,
        64'hffb06ed6_fe0855fe,
        64'h004dbf6a_01f42c5f,
        64'hff621215_0095418f,
        64'hffcf5d8d_fe4e75c0,
        64'h00879438_fff1ddd6,
        64'h0048ad6e_fee423c6,
        64'hffa9bee6_01ebf0d5,
        64'hff2d2a10_007ac11d,
        64'hff241277_fe8bd879,
        64'h00d0c68a_00c583fa,
        64'h00b24f0e_ffe88782,
        64'h0064ff77_feaa7e48,
        64'hff445b7c_ff3895fc,
        64'hffee0cdf_01b1d7d7,
        64'hff328a02_ff82831f,
        64'hfffb33f0_017d1fc9,
        64'h00e2fe54_000a88fa,
        64'hfff50dd9_ffdb623c,
        64'hff9176be_01ae4589,
        64'hff3d85d0_fea365e2,
        64'hff377f26_008f1970,
        64'hff3135bd_ff347e16,
        64'hff0116db_017041b6,
        64'hffba15e4_fefe5831,
        64'hff12f676_00233c86,
        64'h0031c612_00f81893,
        64'h0008450c_fe9c2b1c,
        64'h0051c1e8_01affed5,
        64'hfff759ff_ff1960e8,
        64'hff557d0a_003cccba,
        64'hff9be6ce_0153b61d,
        64'h0001cc7f_ffc78f8a,
        64'hff439371_fe5fafd9,
        64'h00c9be95_0147a1e8,
        64'h00f9d9c7_01e21d48,
        64'h008f0712_ff3b50d6,
        64'hffc6be9a_019b1115,
        64'h00bc6ea6_01078ac2,
        64'hffe47f22_008c4254,
        64'hff34f860_ffa20027,
        64'hff5d7b5a_ff01b443,
        64'hfff8b839_0050b5cd,
        64'hff211717_00e1b7db,
        64'hffb23ee7_00ae5c97,
        64'h00710397_01bbd9c3,
        64'hffbdd2f1_013c1444,
        64'h008df9f7_ffe00546,
        64'hff727e0a_0110875c,
        64'hffa0da25_ff7b4c0f,
        64'h00a531b0_00fad3fd,
        64'hff8ad0d4_ff460efb,
        64'h006468ac_ff74277f,
        64'hff1a55fd_ff17ed0e,
        64'hff57e0ac_fef41f97,
        64'h006ac722_01640ad5,
        64'h0035fbfa_01c136b0,
        64'h003586e4_ff78b2ab,
        64'h00f898d9_ff73c60f,
        64'h006a5cc0_ff174ddf,
        64'hffb9cbba_ff7d5a61,
        64'h008ef586_ffb28c85,
        64'hff05ac54_01ab706a,
        64'h003aa261_010aafe1,
        64'h00e2a7f9_ffb349eb,
        64'hff237ddf_01926540,
        64'hff00d603_01d94513,
        64'hff30c0fd_ff07ff01,
        64'hff42ecc1_001effb3,
        64'hff78f815_013a8f36,
        64'h0011736d_0181cfdb,
        64'h00cd3443_feba914e,
        64'hffaca45b_0005448c,
        64'h0038f1ed_0192c619,
        64'h002a9620_feb63999,
        64'h00fd65da_006671bb,
        64'h00f4b831_ff0d0cec,
        64'h003fa61e_ff824cde,
        64'h008e4f30_fe594a0a,
        64'hfff5cd32_00bb8eec,
        64'hff6692d0_ff2d2ade,
        64'hff166d04_003be0a1,
        64'h008b7f36_01cbfe9e,
        64'h00d39596_fe6008a3,
        64'hff4dde49_01d1f41a,
        64'h0033f4dc_00b180cd,
        64'hffad45ea_ff51b13b,
        64'hff76795d_fead85b7,
        64'hff3e483b_00c54144,
        64'hff728f2f_fff549d2,
        64'h00825355_0173e8e7,
        64'h007f1f23_fee01e24,
        64'h00e2b066_017edc5f,
        64'h00f09d5a_00d34f5e,
        64'h00596162_001b5ad7,
        64'hff278ea2_005ce609,
        64'h0022f5d5_01a70bc0,
        64'h00bc49d0_ff159647,
        64'h007b5524_00600f07,
        64'h006fac70_01185e6e,
        64'hff06d93b_01797141,
        64'h00324e2b_fec10c85,
        64'hffdb0bb1_0070a31f,
        64'h006087b4_01e1cf92,
        64'hfffc921d_fe0016b4,
        64'h00dbdaa5_00510709,
        64'h0073a228_ff0be12a,
        64'h00c3c995_ffcd69b1,
        64'h005cfdd8_0127de44,
        64'hff3fa0c2_00201169,
        64'h002e7a70_ff74da6b,
        64'hff855484_ffbf6363,
        64'hfffe6152_018c05bd,
        64'hff501446_fe441855,
        64'h005dda0d_ff937fa3,
        64'h009f1dd5_01df78f0,
        64'hfff1d176_fecd30d1,
        64'h009a565f_feebe8c3,
        64'h006ab761_ffd58d3d,
        64'hffda03f0_fef543ce,
        64'hff0193c6_01992858,
        64'h00e34a11_ff5ed413,
        64'hff5cb0a5_005492c3,
        64'h007fbff7_00ecdae7,
        64'hff27daf7_003e8962,
        64'hff36abe9_ff7bd734,
        64'h00439303_fe702466,
        64'h009ce60c_008da2d6,
        64'h007cd18a_012a2daa,
        64'hfffdbbd2_ff53630d,
        64'hffab2ec8_ff59b242,
        64'h00c62698_fe849aa7,
        64'hff0a2f44_fed61d0d,
        64'hffea7538_0060da7e,
        64'hff68c678_feb854f5,
        64'h0084a412_0017bb95,
        64'hff908b1b_0126042a,
        64'h00d64f2a_0048190d,
        64'hff489512_fef64331,
        64'h000bda19_ff36b802,
        64'hffd0d599_01533362,
        64'hff21061a_ff60cc93,
        64'hfff33742_004387a0,
        64'h0060f740_014e56ae,
        64'h001c0c18_ff434161,
        64'hff20d68c_ff4c6332,
        64'h00a5f61b_fe7b377b,
        64'hff65d50d_01e87b76,
        64'hff51bed1_0117de0e,
        64'hff03762d_fe19b1a3,
        64'h0026ab9d_ffe2df5e,
        64'hffc79a8a_fe6b2814,
        64'hff3e7346_016dcd8d,
        64'h009af019_ff0e9b21,
        64'h001c3059_ff1e068a,
        64'h00d15488_00b579b0,
        64'hff17717d_ffc290a7,
        64'hfff5fef4_fefe2007,
        64'h00467634_01cba5b0,
        64'hff3a641a_ff149708,
        64'h0057d944_015f101a,
        64'h00640928_00d71fe0,
        64'h00b78975_00ba6346,
        64'hff7c2deb_ff68aaf4,
        64'h008f5cb3_fea93c87,
        64'h00ba09e4_01d06dcf,
        64'h00eda86a_fe205275,
        64'hff32eb4a_ff9663ab,
        64'h002112f8_fee2adf4,
        64'hfff4ed2a_ffe1b464,
        64'hffaf70e3_007dba0f,
        64'hff362587_00ae7452,
        64'hff143607_00e906fc,
        64'hff407aef_00195a9d,
        64'h00660189_fe662adf,
        64'h005b6237_fe24ada9,
        64'hffc0457b_fe86c21f,
        64'h00ccbcd6_0114f8fc,
        64'hffda753c_00c7e2e6,
        64'h00aee24b_01a8de6c,
        64'hff7ebe3e_fea66063,
        64'hff0234db_0163727f,
        64'h00ef0620_ffa47eba,
        64'hff1b1c2d_fe5d3b97,
        64'h009c16d5_fe38ea41,
        64'hff421975_fec2a7e5,
        64'hff134abc_fed7521e,
        64'hff767f45_01f8de7f,
        64'h00928245_fe46487a,
        64'hff115e65_0076b887,
        64'h00f8efeb_fe94ca90,
        64'h00447da5_ffae5089,
        64'h008be584_fec6faba,
        64'h00e9797c_ff132316,
        64'h0014af95_fe99699d,
        64'hffca88ec_fef89840,
        64'h009a4550_fed6fe4b,
        64'h00e9dd63_fe4c86cb,
        64'h0088e4f9_febb3ab6,
        64'h00683a5b_fec840a2,
        64'h0045e79e_012ca8c3,
        64'h00856ed5_ffd003d6,
        64'hff420854_ffa574bd,
        64'h00357f7a_0148eed7,
        64'hffda5392_008c01be,
        64'hff7d8006_ff00ff45,
        64'hffd62aa6_01c94c9f,
        64'h004fd05b_00d64762,
        64'h00dcaaa8_fea45830,
        64'hff242490_ff8fa701,
        64'hff152a82_00e2ac0b,
        64'h008da290_fe9ef8cb,
        64'hff05c693_0138598d,
        64'hff568c82_ffb25cc4,
        64'hffbdf37c_fee44b3b,
        64'hfff1a52a_01282840,
        64'h00a7f767_fe6efdbf,
        64'h008be600_00ab19ce,
        64'h004e4083_00d49e97,
        64'h001cfe83_013440cd,
        64'h00b5092e_00177ce5,
        64'h00e27e34_fe3193dd,
        64'h005c4b5d_ff46888a,
        64'hff08141d_008dc74a,
        64'hff597baa_fef650de,
        64'hff515ce1_fe7394f6,
        64'hff4d05f7_ffe7e29c,
        64'hff971885_fe72c35f,
        64'h0029d879_00844a16,
        64'h00a6f200_fe91b7f4,
        64'hff0eff01_ff253a33,
        64'h00d2ab00_fe097bf4,
        64'h00e7c994_ffd41501,
        64'hff63dce6_00048c98,
        64'h003e3e8a_fe182614,
        64'hff48d9d4_ff2499ec,
        64'h00766691_01b5b5fd,
        64'h007fc5df_00ea16df,
        64'hff7a37d4_ff8010ce,
        64'h0058e45e_fe262868,
        64'hff1efdcf_00a8a968,
        64'h0090cb23_fe7084fa,
        64'h001dc328_fe824e1b,
        64'hff3f3016_fe7fe03b,
        64'hffaa15fe_017f3f10,
        64'h00fe3141_01b7a77f,
        64'h00305cb7_ff447ecb,
        64'h00e909d9_fe32ac19,
        64'h00dbaaf7_01dd4cbf,
        64'hffae20ab_01bac0b7,
        64'hff35cf0b_00b8ee0e,
        64'hff8e034c_009fe18b,
        64'h002f0f42_00194a32,
        64'hffb5624b_01a6a609,
        64'h00ee2f9c_00950026,
        64'hff76a155_00796b8c,
        64'h000111a3_009d9fc8,
        64'hff761037_fff6c6f6,
        64'h00f1765a_fe011ba2,
        64'hfff3d980_fe080d82,
        64'hfff314f1_ff113352,
        64'hff403eb0_fe7731cd,
        64'h008772e3_fe606a83,
        64'hff02505a_ffd7457a,
        64'h00ab419e_ffe925ad,
        64'h0008ae2c_fef57a2d,
        64'h00ec33d3_fe465030,
        64'h00a0e322_0063bdc1,
        64'hff287b32_01080975,
        64'hff6e6000_00aa11a9,
        64'hff95d202_ff6dc17c,
        64'h006916f6_0087fab6,
        64'h00fbc095_ffb2b2ce,
        64'hff1feaeb_009c4e9a,
        64'hff6025d9_010b64b4,
        64'h00c1e6bf_007a74cd,
        64'hff73581a_00acf4f3,
        64'hfff35a09_ff53cffe,
        64'h006cdec5_0125105a,
        64'hffe41170_001c70d4,
        64'hffcea8f7_fe2c0eda,
        64'h00836d9c_0178b265,
        64'h00808d2a_ff789ece,
        64'hff9e0fe3_009f96a6,
        64'h00ce0f7d_005f80be,
        64'hff575d5f_ff8aec27,
        64'hffa1d5aa_fe0dac5f,
        64'h00e97db5_011b0af9,
        64'hffcf874e_0073be0f,
        64'hff330f9b_01bfc19e,
        64'h005e8b46_ff5650ed,
        64'hff6da7df_ff85c5e8,
        64'h00760565_fed60bd4,
        64'hff18dbd7_006f2322,
        64'hffd1bc7e_fea08867,
        64'h001bb52e_0155810a,
        64'hffd29100_01a308fd,
        64'hff0a3459_fe3a0e39,
        64'h005a80ff_01a8e79f,
        64'hff0b8fd4_016da342,
        64'hffb77871_01e41b49,
        64'h001d69a6_fe0c0b9f,
        64'h0059867e_fedb57a2,
        64'h0048adf7_01a2e97b,
        64'hffc9d4b8_0017c01f,
        64'h0041fb18_01944c5e,
        64'h00924832_00951491,
        64'hff17f9c4_ff505243,
        64'h000d9d19_0019c8db,
        64'h0046f228_ff6bf902,
        64'h00d5b96b_01a20587,
        64'h000bd4da_0161494b,
        64'hff1baf89_ff09e5f0,
        64'hffe80f28_fe9633e8,
        64'h000f9bbc_0027fa98,
        64'hff8b603f_ff841b34,
        64'hff5076e2_ff4e89a0,
        64'h00548aa9_ff178d90,
        64'h0088aff1_01f8dc52,
        64'hffa06ba5_fe777edc,
        64'h0004dea0_ffa6b16c,
        64'h00d278c7_fe2d2638,
        64'hff8490d9_ff41f08b,
        64'h00223f94_feb8c225,
        64'h006250c8_0141a0d1,
        64'hffdf74e7_0130fe45,
        64'h00ce1095_fe4b107b,
        64'h00c459f2_feb83be0,
        64'hffc43c7b_fe740dc8,
        64'h0041d91d_fe70db1f,
        64'h00f30e3c_feb9fea3,
        64'hff9bd17f_ff4f80c6,
        64'h006b2586_01ff649a,
        64'h00cf709e_fee0e089,
        64'hff80f7c4_016f2f8a,
        64'h0043403a_0153c4ca,
        64'h004bcea7_017572af,
        64'h00cc6862_01219972,
        64'hff4eda0d_01e18d8f,
        64'h00a283b4_ffd6b26e,
        64'hff8fcea6_01e11b10,
        64'hff766194_013a2fa7,
        64'h008ce74d_fe0766e7,
        64'hff874446_ffea48b9,
        64'h001d5e27_ff88ea86,
        64'h006f4d4c_ff2ec618,
        64'h004c24fc_005959b2,
        64'hffdc6d01_fe2c1e1c,
        64'h004a5ff5_00e07c43,
        64'hffa8fdd6_fe998651,
        64'hff06ef09_015e2f03,
        64'hff70fef2_001379fa,
        64'h00e5f2ea_00862460,
        64'h006ebaa4_01075817,
        64'h0025a4a8_0062c526,
        64'hff200be0_0000dfaa,
        64'h009fdac2_00039d51,
        64'hff419eb3_feb6ccdd,
        64'h00befc36_01ffa7b3,
        64'h00e61d6e_00d73e9d,
        64'h007e1b13_ff144b16,
        64'h00c763db_00df182b,
        64'h00807ccc_0139e457,
        64'h000d1a49_fe934017,
        64'h000f26dc_ff8f10b5,
        64'h0005769f_00801406,
        64'hff10c729_0196cf14,
        64'hff7981ed_fe518a43,
        64'h00f218da_ff8a20bc,
        64'h00cff668_004341ba,
        64'hfffa064d_0080e149,
        64'hff48acb8_ffc0c753,
        64'h00929db7_00ea8aeb,
        64'h007dc000_0092b281,
        64'h00e2ef78_ff9fc040,
        64'h006491dc_01f9972d,
        64'hff601648_00c47c89,
        64'h00bc4bfc_ff4cc5ac,
        64'hffbaaaa8_01778b0f,
        64'h001de61b_fe19a95e,
        64'h00f3af1a_012c477d,
        64'h007fb1bc_00e7f04c,
        64'hff6d8171_0047f033,
        64'hff047609_fec4d7a3,
        64'h001c3111_01c0dde3,
        64'hffaee50b_ffb406ee,
        64'hff84d2e5_fe5112f4,
        64'hff494867_fe473905,
        64'h00f0ba64_fffeed25,
        64'h0047b37f_01f3bc04,
        64'h00a523ff_fedef7a4,
        64'hffcbd1bd_00dafee2,
        64'h00a4f871_00e6c4a3,
        64'hffc75369_0012331a,
        64'h00fdea2f_01214193,
        64'h00117e07_fe599b1c,
        64'hff4f799b_fea91948,
        64'hffa651a3_ffdbd96c,
        64'hff75e632_001ebb93,
        64'hff7ef7f9_00c1ec05,
        64'hff867863_ff0f2f22,
        64'hffc61d5f_ff53a490,
        64'h00587498_ffa963ea,
        64'h0071a0ae_0085955d,
        64'hff5459c5_ff0fffec,
        64'hff983760_0116fbe9,
        64'h003b81d5_fecfce4e,
        64'h00b00fd5_fe56c2b0,
        64'h007b3b75_014cf572,
        64'hffd907a0_feded49c,
        64'h0076140a_0073a463,
        64'h00a315c1_0078433c,
        64'hffd0372a_fed58f0e,
        64'h001a4304_01b03bce,
        64'hffd54770_0013b087,
        64'h00b108cb_fe5dc12c,
        64'h007d19f2_feca62d1,
        64'h004ce9e0_0007380b,
        64'hffb06cd7_005b3728,
        64'hffc07236_01fdad52,
        64'hff2b19ae_00302ff3,
        64'h00b4654a_00b24cc2,
        64'hff6edf6c_01230680,
        64'hff0593a4_ff1ed457,
        64'hffa3d763_ff193227,
        64'hff15ee6f_ffb930b9,
        64'hff24c845_01e7793d,
        64'hff6f5d15_00308304,
        64'hffb99ef9_01a37d0b,
        64'h00c035cf_ff179b23,
        64'h007cc123_01f1b929,
        64'h00cb4d62_ff4ec565,
        64'h00100fb4_01d0ca68,
        64'hffc5344f_00ec3269,
        64'h0007e3a0_00ca15f1,
        64'hff652a7f_ff124933,
        64'hffddff4f_fe2dcc7f,
        64'hffcc2e65_010f7059,
        64'h00ba6c81_01260b31,
        64'hffcbf45a_01588770,
        64'h003bd659_017be2cf,
        64'hff09e2e1_01eaec41,
        64'h0082627a_009fe274,
        64'h0058d3e0_018d300c,
        64'h00acf6d1_01c95045,
        64'h0007020c_016a2e51,
        64'h0034751f_001764b6,
        64'hff5812a2_fedcbfa7,
        64'hffce9258_014a6098,
        64'h007c0d1d_ff710376,
        64'hff85e324_fe7d6613,
        64'hff268423_fe5bcfe7,
        64'h001a869b_00288675,
        64'h002b7234_01a97b29,
        64'hff5763ec_fe29361b,
        64'hff662c42_00e822ac,
        64'hff58a308_fe9c572e,
        64'hff27d7ef_ffa496cc,
        64'hffd7e7b0_ff55f38d,
        64'hff0baa25_ff85894f,
        64'hffa308b5_010c3a46,
        64'h00840b4f_feeb9302,
        64'h00f780bb_007ca8f8,
        64'hff796e4e_0019e04f,
        64'h00f01c88_0165e545,
        64'h00f55f9f_01914626,
        64'hffc34720_00b49bfa,
        64'hff226d3e_00670301,
        64'h00516c21_00089b61,
        64'h009f05ee_ff919798,
        64'hffd50c63_0083d337,
        64'h006cdc68_ff18b570,
        64'hff646d9f_019bffed,
        64'hff170d2c_ff14832c,
        64'h00aa2b8f_004bbfe6,
        64'h0026697c_ff981e32,
        64'h00291d28_00846a89,
        64'h00b218ec_000afaf5,
        64'h007ab299_01b080fd,
        64'h0052b667_fe87e831,
        64'hff9cc51a_ff56ae56,
        64'h00afd784_0124422a,
        64'h000596d7_fe48efca,
        64'h00902ca5_fe609520,
        64'h009e2af5_0086a2db,
        64'h00486722_01e6b024,
        64'h005381b7_ff096ab8,
        64'hff041374_002fe9c6,
        64'h00ef6722_00a94891,
        64'hff9d3c53_fe308652,
        64'h00e10148_01931635,
        64'h009a07e3_00933979,
        64'h00ffcbe8_01ebd5dc,
        64'hff7a8b94_00de1545,
        64'hff611854_011a6613,
        64'hfff7b420_015528d5,
        64'hff24bd9e_0134f027,
        64'h009e3faf_fed4eaea,
        64'h003733fa_0085b6b5,
        64'hff60a88d_015b0d17,
        64'hffdc479a_010ffc4b,
        64'hffcbdf67_fee4756d,
        64'h005233d6_00d34c9f,
        64'hff900e3e_fe310813,
        64'h00bb8158_fe74f9d2,
        64'h00d48aa3_01e787fb,
        64'h00b40524_fef0d6e0,
        64'h004e055e_fe297912,
        64'h00b84793_00cbaec9,
        64'h00e187cb_fe005845,
        64'h00e30859_ffd59eba,
        64'h00957928_fe7dd6b7,
        64'hfff51f1b_fe2cfb89,
        64'h00061421_ff2f0ef2,
        64'hff052b75_ff971be9,
        64'h00cb1ce2_00dae87f,
        64'h009e51e1_001e752b,
        64'h00fb9cc0_00f2685d,
        64'h008c81ac_00d6f10d,
        64'hffd59e3c_01cdaeb9,
        64'hffd2deea_004c0660,
        64'h006d6653_ffbc8989,
        64'hff3adca3_0012fcdc,
        64'hffbeef87_01450c51,
        64'hff3b603e_0075236b,
        64'h00a0ada9_0164a81d,
        64'h001f511d_004346d1,
        64'h002a1c78_0070c6aa,
        64'hffc3bb5c_0164861b,
        64'hff4afae7_01922275,
        64'hffe8542e_fe990fc4,
        64'h00d3165f_006691ae,
        64'hff06ee22_ffb726d1,
        64'h00427eec_00587c8f,
        64'h0006d93a_ff383dea,
        64'hffe12315_ff368116,
        64'h006dd523_001af903,
        64'hff2406aa_ff183c51,
        64'h003e6049_fe0e2d44,
        64'h007fd0d2_0087f2bb,
        64'hff118d6c_feefcc8a,
        64'hff562992_01fe1e57,
        64'hff04dde4_0166feac,
        64'hff214d99_00033f41,
        64'h000c214d_00ac083a,
        64'hffa49ec7_ffc147be,
        64'h00b4a771_00244e58,
        64'h003f3b04_00f01e02,
        64'h002a2c35_00045af7,
        64'h00ff6b67_ff048d48,
        64'hff8df725_ff9323eb,
        64'h00bd812c_fea6ae05,
        64'hffd26ddc_ff96fb12,
        64'h000dfa41_fe393100,
        64'hff28c561_01cee60a,
        64'hff5d6f9b_ff7dae3e,
        64'h003ef126_fefce360,
        64'hffbdfa4f_0020796c,
        64'h00f71188_004ee03b,
        64'hff1c8bc3_012d9b4d,
        64'hff1a825c_01227be5,
        64'h00df09ab_016f1ea5,
        64'h004ad7f9_fefa048f,
        64'hffb6d55b_ffe8fcd0,
        64'h0091f285_00777a1f,
        64'h00d5a4ba_ff0b078d,
        64'h0048cb66_fe3ddb34,
        64'h00fe802a_ffe71383,
        64'hff9dba8c_00c34460,
        64'hffe107cf_fe3e639d,
        64'h00e07efb_ff4cca28,
        64'hfffb82c3_fe9d5294,
        64'h00005d4f_019f7cd7,
        64'hff98895f_00112680,
        64'h00ac824b_ffa3e253,
        64'hff8cb03d_ff59d623,
        64'hff19c81e_ff2f5ee4,
        64'h00094874_ff67a636,
        64'hff4acdea_016bdc4d,
        64'h00a29a50_00190280,
        64'hffbdd61d_00efc1f5,
        64'hffde3c78_01415b8a,
        64'h007efa96_fec3b190,
        64'hff33286c_01f8290b,
        64'hfff03baf_fecc1c5a,
        64'hff7cb7a7_fe04e5f7,
        64'h00a67f50_00d1add9,
        64'hffafd641_01730908,
        64'hff9193c7_000a0645,
        64'hff10bc61_ffbc4851,
        64'h0000b60b_fea6ac68,
        64'h002572c5_002465a3,
        64'h00dcdd9d_0075c652,
        64'hffe08675_fe5e41d5,
        64'hffbe8195_00d2558e,
        64'h006769da_fe19e497,
        64'h002ceb95_feafdedd,
        64'h00bf671c_01e5f758,
        64'h002e73c2_fe2eb09e,
        64'h0085e88b_01b1d139,
        64'hff855276_feb4ffe8,
        64'h00dee126_ffdd95c2,
        64'h0017f0ef_004535d8,
        64'hff6fd7ed_feab6767,
        64'h001d4f81_ff995b77,
        64'hffca0524_fefc643d,
        64'hffc2cbd4_fe71ecb8,
        64'h00520a74_fea83fc5,
        64'h004d85f8_01f95b3e,
        64'hff61131e_0164f97a,
        64'h00264e40_000ae79b,
        64'hffd1859a_0185f7d4,
        64'h00ce5d6f_00a5ecc3,
        64'h00bb2397_fef607c0,
        64'hff7fd2dc_fef2395b,
        64'h00ad44de_008a22c7,
        64'hffe927e7_00c10834,
        64'h0053ee98_ff34793b,
        64'h00454d01_0171203a,
        64'hff1aee58_01b19045,
        64'hff5798b3_00f87421,
        64'hff50a172_fe5a2fd0,
        64'hff59b5e2_fe34586e,
        64'h00459417_ff1ef6e6,
        64'h001268f5_01bd61d0,
        64'hff65a2cc_fe8fc7e2,
        64'h00f84a33_00586617,
        64'h00979873_febed670,
        64'hffc121c0_006fe423,
        64'h00304590_0099753f,
        64'hff68cd6c_ffd44c92,
        64'h00f109df_01be5fde,
        64'h000efe6f_fef55080,
        64'h00ddee8d_fe69d31e,
        64'hff11eddc_01a8f52c,
        64'hff1bd102_0048e195,
        64'hff8aa821_ff58c805,
        64'h00431a5c_0112e865,
        64'hff76168e_01cf5235,
        64'hff4d3f27_ffed4f5a,
        64'h0004946c_ffed2d89,
        64'hff1105c8_0106e4c7,
        64'h00c35db6_fef03d31,
        64'h00b730a2_fe0ff4ae,
        64'hff42d1c5_fea19712,
        64'h00f85e34_00475dab,
        64'h00d8d512_01aa515e,
        64'hffb74df5_009a00ef,
        64'hffe72a5c_ffdbb5d4,
        64'h00637a58_014742da,
        64'h00b3b44a_fe22a5da,
        64'hff374399_ff2f9c30,
        64'h009a41f1_01c2ecc5,
        64'hffd2ac6d_fe090c87,
        64'h00b62a33_fee28dc6,
        64'hffc45e65_00fafcf8,
        64'h007d7672_01a2911a,
        64'h00ea4093_fe1320e0,
        64'h00386585_ffa0d637,
        64'h003c23fc_fe58f5da,
        64'h00070dab_ff1f3c55,
        64'hffd77b7d_ff9234d9,
        64'h0024579e_fe061bce,
        64'h00a5f626_01ce332f,
        64'h00d9c323_01b2cc0e,
        64'hffbf1444_fe058b37,
        64'hffd65981_00dd3e8f,
        64'hffea7eec_01c6a0f9,
        64'h0014ea54_fe20dd2c,
        64'h0077adf4_fecc0d7d,
        64'h003829f5_00935e30,
        64'h00db7200_01b8b3b5,
        64'h0075bb75_01d2e531,
        64'h00fc13bd_013b27c9,
        64'h00192c3a_01b28085,
        64'h0099ddd1_0074f74e,
        64'hffcb26ab_fe3221b1,
        64'hff186faa_fe9283c9,
        64'h004fce36_01294114,
        64'h00542e49_01d1c0d5,
        64'hffd59cee_001a4d63,
        64'h00973425_004ea3d2,
        64'h0042e3a4_01a9f0d6,
        64'h003c6a7d_fe512584,
        64'h003bc145_fef9c380,
        64'h001a0d0e_ff6030b6,
        64'hff0c99c1_feea4b71,
        64'h00e2d931_001ae418,
        64'hff109761_002e7390,
        64'h004553b9_015d6f8a,
        64'h00213e91_00e72933,
        64'h0001ad9f_ff7d8ca4,
        64'hff4795ef_ff6a2cc4,
        64'hff17b00d_fedb346d,
        64'h0059a737_fe6c9c56,
        64'h00480645_01f10742,
        64'hff3bbade_ff157144,
        64'hff0eaafa_fe96b3bb,
        64'h00d35683_01b3858e,
        64'hffbda72d_009c3820,
        64'h003e85ef_fe3f9797,
        64'h00f6fc60_012a8298,
        64'h005529fa_ff3eb1b5,
        64'h00be7c68_fe788e5c,
        64'h0064a088_ff540053,
        64'h008a5939_0136eff2,
        64'h0060b0e9_0047d6ba,
        64'h00a51734_ff146e20,
        64'h00dd7ba3_01f5862d,
        64'h00bfec45_fe354123,
        64'h001e3af7_01a05442,
        64'h00af1102_00a5bb33,
        64'hfffe7433_fff63554,
        64'hffc56bbb_01ee7c88,
        64'h002b4494_01ba78e5,
        64'h002bdae6_002e4b42,
        64'h00fefa71_0076ff1c,
        64'h009e4cfd_00c7445a,
        64'h0093587d_0071e683,
        64'h00a05073_00c9fa26,
        64'hff8ab308_ff5532c0,
        64'hff814281_016818bf,
        64'hffa03a44_00321e58,
        64'h00e4f947_fe469efe,
        64'hff0a9265_019d971c,
        64'hffa3efe9_00a7050e,
        64'h00d46e64_fefc09b2,
        64'hff68a09b_fef12b9b,
        64'h0098da2e_0072a2c6,
        64'h00f2db4c_0162508d,
        64'hff10e1af_ff4c4296,
        64'hffa4cfc3_01d0d89c,
        64'h00aae456_007555be,
        64'hff4c5026_00f98d11,
        64'hff4bd6bd_00ef4d50,
        64'hffef2e0e_ff4faacc,
        64'h0047fa29_00fcd265,
        64'hffe85938_01b9a810,
        64'hff1e9823_01a80150,
        64'hff016732_00096a11,
        64'hff874432_017155e5,
        64'hff6c2a13_00ee9743,
        64'hffc06bd7_ff13ea51,
        64'hff6e6a02_ffd04206,
        64'hff3d6a31_00db05af,
        64'h00eaecd6_01ef087f,
        64'h00aa2ce9_019b7a72,
        64'hffaed657_fe669c92,
        64'h00aabc14_ff11b5d9,
        64'hff6e37ab_fe3cae04,
        64'h00627305_019ed153,
        64'h00695811_feb4d5bb,
        64'hff643019_fffa87d3,
        64'hffc5cb55_ff4d32f1,
        64'hffd60703_fe7d1a76,
        64'h00b3d080_feb6b245,
        64'hff39ff25_ff3c71ea,
        64'hffbc45ee_fe89f0c6,
        64'h00b50b43_01bee5ef,
        64'hff43598c_009b67a1,
        64'hff1e6556_0093d579,
        64'h00448162_ff7aaa7b,
        64'hff13f4be_01298f81,
        64'h004cf4b8_00c21a34,
        64'h008f8a0a_fff4e67c,
        64'h002e8a06_ffd673a2,
        64'h000e4176_ff409151,
        64'h001f3e75_ffa33d4c,
        64'hff4ca4e1_01a44c32,
        64'h003d42c3_ff3e4cb7,
        64'h0037dc60_01c325f8,
        64'hff24f1bd_018c3b85,
        64'hff447585_fe10ae4e,
        64'hff084066_ff2d3eca,
        64'hffd64271_fface2bd,
        64'h0071b9ff_ffddcbb3,
        64'h009d8be7_ffd0b529,
        64'hff0ed735_00218d06,
        64'hffd7eea1_00180404,
        64'hffb25193_ff4e0a6f,
        64'hff2154c9_fe1ac081,
        64'h00f36192_fe8ccf1e,
        64'hff8788a4_017f12de,
        64'h00e565b8_fedefd61,
        64'hfff2d4d1_fe19230a,
        64'h0068c4e1_008da49a,
        64'hffb300c5_ffcfeab3,
        64'hff25ee9c_ffdaa098,
        64'hff0c745e_ff9bfc49,
        64'hffa7e533_0090df9b,
        64'hff8efc6f_fe8e2a6c,
        64'h0028465d_ff2ea38b,
        64'h00099e21_fed17602,
        64'h0094f3a2_01591955,
        64'h00ad5969_febbf3af,
        64'h004cdbbb_01ed6a0e,
        64'hffc04ecd_fe7fbf93,
        64'h008d3f60_feec346f,
        64'h00482a6f_0107097e,
        64'hff07ba08_fefe12ce,
        64'h00d5ade7_ffdb77ee,
        64'h003088a9_fe007f6d,
        64'h00f71955_fe2b53e0,
        64'hff290886_0088ccdb,
        64'hff1a8622_000c7ad3,
        64'hff099417_00949b05,
        64'h00cb317f_016089e9,
        64'h0062ad66_00029d5c,
        64'h00eff474_003aaab5,
        64'h008deb95_00fb5ace,
        64'hff4bb844_0070262c,
        64'hffd6c092_01864348,
        64'hff09d6ac_fe2546d9,
        64'hfff5e228_ff42388c,
        64'hff703407_ff9767fb,
        64'h00781181_01c4e5f8,
        64'hffc02123_fe802af1,
        64'hffcf05c8_0021b009,
        64'hff60d55f_ff7e14ca,
        64'hffd4cf17_ff8bfe10,
        64'hff4538cf_fe45e0d7,
        64'hff3a2fe4_0045af2e,
        64'hff270169_011fadca,
        64'hff91f2d9_01e30474,
        64'hff5eb045_fe628207,
        64'hffb7a902_00337e6e,
        64'hff885f81_ff9d8077,
        64'h00d2e7b5_ff38add8,
        64'hffeb39d6_0119e4e3,
        64'h0086f5b6_fe99427a,
        64'hff7a8de2_00d8b366,
        64'hff99e2aa_fea8632f,
        64'hffea7eec_01c6a0f9,
        64'h0014ea54_fe20dd2c,
        64'h0077adf4_fecc0d7d,
        64'h003829f5_00935e30,
        64'h00db7200_01b8b3b5,
        64'h0075bb75_01d2e531,
        64'h00fc13bd_013b27c9,
        64'h00192c3a_01b28085,
        64'h0099ddd1_0074f74e,
        64'hffcb26ab_fe3221b1,
        64'hff186faa_fe9283c9,
        64'h004fce36_01294114,
        64'h00542e49_01d1c0d5,
        64'hffd59cee_001a4d63,
        64'h00973425_004ea3d2,
        64'hff0eaafa_fe96b3bb,
        64'h00d35683_01b3858e,
        64'hffbda72d_009c3820,
        64'h003e85ef_fe3f9797,
        64'h00f6fc60_012a8298,
        64'h005529fa_ff3eb1b5,
        64'h00be7c68_fe788e5c,
        64'h0064a088_ff540053,
        64'h008a5939_0136eff2,
        64'h0060b0e9_0047d6ba,
        64'h00a51734_ff146e20,
        64'h00dd7ba3_01f5862d,
        64'h00bfec45_fe354123,
        64'h001e3af7_01a05442,
        64'h00af1102_00a5bb33,
        64'hff68a09b_fef12b9b,
        64'h0098da2e_0072a2c6,
        64'h00f2db4c_0162508d,
        64'hff10e1af_ff4c4296,
        64'hffa4cfc3_01d0d89c,
        64'h00aae456_007555be,
        64'hff4c5026_00f98d11,
        64'hff4bd6bd_00ef4d50,
        64'hffef2e0e_ff4faacc,
        64'h0047fa29_00fcd265,
        64'hffe85938_01b9a810,
        64'hff1e9823_01a80150,
        64'hff016732_00096a11,
        64'hff874432_017155e5,
        64'hff6c2a13_00ee9743,
        64'hffbc45ee_fe89f0c6,
        64'h00b50b43_01bee5ef,
        64'hff43598c_009b67a1,
        64'hff1e6556_0093d579,
        64'h00448162_ff7aaa7b,
        64'hff13f4be_01298f81,
        64'h004cf4b8_00c21a34,
        64'h008f8a0a_fff4e67c,
        64'h002e8a06_ffd673a2,
        64'h000e4176_ff409151,
        64'h001f3e75_ffa33d4c,
        64'hff4ca4e1_01a44c32,
        64'h003d42c3_ff3e4cb7,
        64'h0037dc60_01c325f8,
        64'hff24f1bd_018c3b85,
        64'h00901b67_01c56e00,
        64'hff9ce332_ff407977,
        64'h00f3d130_00038052,
        64'h00d4141e_fe2add7b,
        64'hffa6e50a_feb2f159,
        64'h00ae0c92_0004fc1e,
        64'hffe1656a_fe804c9f,
        64'hfffbd7a7_00bd0c60,
        64'h0035697f_008f189e,
        64'hff86c9d3_fe0ea0b0,
        64'hff480db4_fee2b700,
        64'hffce7199_ffa03cbc,
        64'hff79e898_0001c029,
        64'h006a0a0f_ff156ebd,
        64'h00d37285_ff5978b6,
        64'h0000f02f_f06f8082,
        64'h61756db2_6d526cf2,
        64'h7c127bb2_7b527af2,
        64'h6a1669b6_695664f6,
        64'h741670b6_7f010113,
        64'hbd79c60f_f0ef8522,
        64'h85da963e_078d8613,
        64'h078e40f6_07b30047,
        64'h961340f0_07bb4017,
        64'hd79b0197_07bb01fc,
        64'hd71bacdf_d0ef1228,
        64'h85a28652_ad7fd0ef,
        64'h020885a6_864aae1f,
        64'hd0ef8562_85d28626,
        64'haebfd0ef_855a85a2,
        64'h864ab5d5_9f7ff0ef,
        64'h852285da_963e1f9c,
        64'h0616963e_00279613,
        64'h40f007bb_4017d79b,
        64'h019707bb_01fcd71b,
        64'hb1bfd0ef_122885a2,
        64'h8652b25f_d0ef0208,
        64'h85a6864a_b2ffd0ef,
        64'h856285d2_8626b39f,
        64'hd0ef855a_85a2864a,
        64'hbf3dc5ef_f0ef8522,
        64'h85da963e_078d8613,
        64'h078e40f6_07b30047,
        64'h9613401c_d793b61f,
        64'hd0ef1228_85a28652,
        64'hb6bfd0ef_020885a6,
        64'h864ab75f_d0ef8562,
        64'h85d28626_b7ffd0ef,
        64'h855a85a2_864af990,
        64'h51e3000a_8c83ae0f,
        64'hf0ef8522_85da963e,
        64'h1f9c0616_963e0027,
        64'h9613401c_d793ba9f,
        64'hd0ef1228_85a28652,
        64'hbb3fd0ef_020885a6,
        64'h864abbdf_d0ef8562,
        64'h85d28626_bc7fd0ef,
        64'h855a85a2_864afb90,
        64'h5fe30009_8c83ef2f,
        64'hf0ef8522_85de153d,
        64'h01631afd_be7fd0ef,
        64'h19fd85a6_864a6522,
        64'hbf3fd0ef_85d28626,
        64'h6502bfdf_d0ef855e,
        64'h85a2864a_100c9b63,
        64'h09904363_000a8c83,
        64'h0c0c9a63_a825028b,
        64'h0c130284_0a130504,
        64'h04930784_09131ef1,
        64'h0d1300e7_8ab31d9c,
        64'h00e789b3_1b9c00c7,
        64'h8b3397da_8e068793,
        64'h7c0b0b13_00c78433,
        64'h081097a2_8e068793,
        64'h720b0413_66857b7d,
        64'hd67517fd_0007c603,
        64'h1cb70263_377dea01,
        64'h16fd0006_c603a801,
        64'h55fd0ff0_07133ef1,
        64'h06932ef1_0793e98f,
        64'hd0efe43e_853e050b,
        64'h8793ea4f_d0efe03e,
        64'h853e028b_8793e86f,
        64'hd0ef855e_c9ffd0ef,
        64'h00278533_865a122c,
        64'h8c8c0793_a15fd0ef,
        64'h020c0027_85338a0c,
        64'h0793c93f_e0ef85ca,
        64'h00278533_8626878c,
        64'h0793f0ef_d0ef85ca,
        64'h86260027_8533850c,
        64'h0793cddf_d0ef1228,
        64'h85a2864e_ce7fd0ef,
        64'h020885d2_8656cf1f,
        64'hd0ef854a_85ce8652,
        64'hcfbfd0ef_852685a2,
        64'h8656c54f_f0ef8522,
        64'h0a8c7b01_0613d11f,
        64'hd0ef122c_865a0027,
        64'h8533828c_0793a87f,
        64'hd0ef020c_00f10533,
        64'h80078793_6785d07f,
        64'he0ef7d81_051385ca,
        64'h8626f7ef_d0ef85ca,
        64'h86267b01_0513d49f,
        64'hd0ef1228_85a2864e,
        64'hd53fd0ef_020885d2,
        64'h8656d5df_d0ef854a,
        64'h85ce8652_d67fd0ef,
        64'h852685a2_8656cc0f,
        64'hf0ef8522_0a8c7101,
        64'h0613d7df_d0ef7881,
        64'h0513122c_865aaeff,
        64'hd0ef7601_0513020c,
        64'hd69fe0ef_73810513,
        64'h85ca8626_fe0fd0ef,
        64'h85ca8626_71010513,
        64'hdabfd0ef_122885a2,
        64'h864edb5f_d0ef0208,
        64'h85d28656_dbffd0ef,
        64'h854a85ce_8652dc9f,
        64'hd0ef8526_85a28656,
        64'hd22ff0ef_85220a8c,
        64'h67010613_ddffd0ef,
        64'h6e810513_122c865a,
        64'hb51fd0ef_6c010513,
        64'h020cdcbf_e0ef6981,
        64'h051385ca_8626843f,
        64'hd0ef85ca_86266701,
        64'h0513e0df_d0ef1228,
        64'h85a2864e_e17fd0ef,
        64'h020885d2_8656e21f,
        64'hd0ef854a_85ce8652,
        64'he2bfd0ef_852685a2,
        64'h8656d84f_f0ef8522,
        64'h0a8c5d01_0613e41f,
        64'hd0ef6481_0513122c,
        64'h865abb3f_d0ef6201,
        64'h0513020c_e2dfe0ef,
        64'h5f810513_85ca8626,
        64'h8a5fd0ef_85ca8626,
        64'h5d010513_e6ffd0ef,
        64'h122885a2_864ee79f,
        64'hd0ef0208_85d28656,
        64'he83fd0ef_854a85ce,
        64'h8652e8df_d0ef8526,
        64'h85a28656_de6ff0ef,
        64'h85220a8c_53010613,
        64'hea3fd0ef_5a810513,
        64'h122c865a_c15fd0ef,
        64'h58010513_020ce8ff,
        64'he0ef5581_051385ca,
        64'h8626907f_d0ef85ca,
        64'h86265301_0513ed1f,
        64'hd0ef1228_85a2864e,
        64'hedbfd0ef_020885d2,
        64'h8656ee5f_d0ef854a,
        64'h85ce8652_eeffd0ef,
        64'h852685a2_8656e48f,
        64'hf0ef8522_0a8c4901,
        64'h0613f05f_d0ef5081,
        64'h0513122c_865ac77f,
        64'hd0ef4e01_0513020c,
        64'hef1fe0ef_4b810513,
        64'h85ca8626_969fd0ef,
        64'h85ca8626_49010513,
        64'hf33fd0ef_122885a2,
        64'h864ef3df_d0ef0208,
        64'h85d28656_f47fd0ef,
        64'h854a85ce_8652f51f,
        64'hd0ef0284_89138526,
        64'h85a28656_00e784b3,
        64'h081897a6_8e0c0793,
        64'h7c048493_ebeff0ef,
        64'h85220a8c_1f90f79f,
        64'hd0ef03a8_85a2864e,
        64'hf83fd0ef_130885d2,
        64'h8656f8df_d0ef1aa8,
        64'h85ce8652_f97fd0ef,
        64'h02840993_05040a13,
        64'h0a8885a2_8656ac3f,
        64'hf0ef0784_0a938522,
        64'h0a8c00e7_84330818,
        64'h97a28e0c_07937204,
        64'h841374fd_6c05d2ff,
        64'hd0ef1308_85cad37f,
        64'hd0ef1aa8_85a6d3ff,
        64'hd0ef0a88_85a2fe1f,
        64'hd0ef4681_05130784,
        64'h0593865a_d55fd0ef,
        64'h050d8b13_58ad8d93,
        64'h44010513_85ca0000,
        64'h0d970504_0913fdff,
        64'he0ef4181_051385a6,
        64'h8622a57f_d0ef1f88,
        64'h85a68622_02840493,
        64'hc54ff0ef_1d8885a6,
        64'hc5cff0ef_843284b6,
        64'h1b888baa_81010113,
        64'hea6aee66_e66ef262,
        64'hf65efa5a_fe56e2d2,
        64'he6ceeaca_eea6f2a2,
        64'hf6867149_80826165,
        64'h7ae26a06_69a66946,
        64'h64e67406_70a6aabf,
        64'hd0ef8556_002c8656,
        64'h848ff0ef_8552002c,
        64'h8656abff_d0ef854e,
        64'h85d2864e_85cff0ef,
        64'h852285d2_864ead3f,
        64'hd0ef0028_85a28622,
        64'h89afe0ef_85220504,
        64'h85930509_06138a8f,
        64'he0ef8556_07890593,
        64'h07848613_07840a93,
        64'h8bafe0ef_854e85ce,
        64'h864a8c4f_e0ef8552,
        64'h85a20289_06130504,
        64'h0a138aaf_f0ef854e,
        64'h85d28626_b21fd0ef,
        64'h02850993_842afc56,
        64'he4cef0a2_f4868626,
        64'h893285d2_e8ca0285,
        64'h8a1384ae_e0d2eca6,
        64'h71598082_22010113,
        64'h6c5e6bfe_7b1e7abe,
        64'h7a5e79fe_20013903,
        64'h20813483_21013403,
        64'h21813083_fb799ee3,
        64'h090992cf_e0ef2989,
        64'h855a1a0c_0ab0938f,
        64'he0ef8552_030c1330,
        64'h942fe0ef_85560aac,
        64'h031094cf_e0ef8526,
        64'h1a0c1330_a71ff0ef,
        64'h1a0885a6_8622e68f,
        64'hf0ef8522_4019d593,
        64'h00090603_04000b93,
        64'h4981974f_e0ef855a,
        64'h1a0c0ab0_97efe0ef,
        64'h8552030c_1330988f,
        64'he0ef8556_0aac0310,
        64'h992fe0ef_85261a0c,
        64'h1330cb7f_f0ef1a08,
        64'h192c9a4f_e0ef0228,
        64'h030c1330_9aefe0ef,
        64'h11880aac_03109b8f,
        64'he0ef1928_1a0c1330,
        64'hcddff0ef_1a08192c,
        64'h9cafe0ef_0228030c,
        64'h13309d4f_e0ef1188,
        64'h0aac0310_9defe0ef,
        64'h19281a0c_1330d03f,
        64'hf0ef1a08_192c9f0f,
        64'he0ef0228_030c1330,
        64'h9fafe0ef_11880aac,
        64'h0310a04f_e0ef1928,
        64'h1a0c1330_d29ff0ef,
        64'h1a08192c_f7dfd0ef,
        64'h022885d2_f85fd0ef,
        64'h118885d6_f8dfd0ef,
        64'h192885a6_fb899de3,
        64'ha32fe0ef_855a1a0c,
        64'h0ab00989_a3efe0ef,
        64'h8552030c_1330a48f,
        64'he0ef8556_0aac0310,
        64'ha52fe0ef_85261a0c,
        64'h1330b77f_f0ef1a08,
        64'h85a68622_f6eff0ef,
        64'h85224015_d59b013b,
        64'h85bb0009_8603413b,
        64'h8bbb0419_0c13c6ff,
        64'hd0ef4b85_00110993,
        64'h855a0784_8b13ca9f,
        64'hd0ef8552_05048a13,
        64'hcb3fd0ef_8556c8ff,
        64'hd0ef02f1_0fa39fb1,
        64'h02848a93_852603f1,
        64'h4783fcd5_1ce3fef6,
        64'h8fa39f8d_0046159b,
        64'h0ff77613_87114187,
        64'h571b0187_171b0087,
        64'h871b0ff7_f7939fb9,
        64'h06850006_c7834701,
        64'h86ca03f9_0513fee4,
        64'h14e3fef7_1f238fd5,
        64'h8bbd0086_969b0047,
        64'hd69b0585_07090005,
        64'hc783874a_008084aa,
        64'hebe2efde_f3daf7d6,
        64'hfbd2ffce_20113c23,
        64'h20913423_20813823,
        64'h890a2121_3023de01,
        64'h01138082_610d64aa,
        64'h644a60ea_00f40fa3,
        64'h8fa90075_151b01f4,
        64'h4783e54f_f0ef1808,
        64'hbccff0ef_852208ac,
        64'hb52fe0ef_08a80284,
        64'h85930030_b5efe0ef,
        64'h180885a6_0030d75f,
        64'he0efed06_05058593,
        64'h002884ae_842ae526,
        64'he9227135_8e4fe06f,
        64'h610564a2_05048593,
        64'h60e26442_05040513,
        64'h8f8fe0ef_02840513,
        64'h02848593_904fe0ef,
        64'h84ae842a_e426e822,
        64'hec061101_baefe06f,
        64'h61050506_061394c6,
        64'h061364a2_07848513,
        64'h00001617_690260e2,
        64'h64420784_0593936f,
        64'he0ef0504_85130504,
        64'h0593bb2f_f0ef0284,
        64'h851385ca_8622e2bf,
        64'hd0ef84aa_e426ec06,
        64'h85ca842e_862ee822,
        64'h02858913_e04a1101,
        64'h8082610d_64aa644a,
        64'h60eaf27f_f0ef8526,
        64'h002c97af_e0ef08a8,
        64'h05040593_984fe0ef,
        64'h18080284_059398ef,
        64'he0ef842e_e922ed06,
        64'h002884aa_e5267135,
        64'he29fd06f_014160a2,
        64'h64020784_0513e61f,
        64'hd0ef0504_0513e69f,
        64'hd0ef0284_0513e47f,
        64'hd0ef842a_e022e406,
        64'h11418082_61657ae2,
        64'h6a0669a6_694664e6,
        64'h740670a6_c4cff0ef,
        64'h855285d2_8626c56f,
        64'hf0ef8522_002c864e,
        64'hc60ff0ef_852685a6,
        64'h8622ed7f_d0ef854e,
        64'h85a68622_ba1fe0ef,
        64'h002885ce_ee9fd0ef,
        64'h854e85ca_86560284,
        64'h099396ef_f0ef8552,
        64'h05090593_07840a13,
        64'hbc5fe0ef_852685d6,
        64'hbcdfe0ef_02890a93,
        64'h05050493_842afc56,
        64'he0d2e4ce_eca6f0a2,
        64'hf486892e_e8ca7159,
        64'hf03fd06f_014160a2,
        64'h64020504_0513f11f,
        64'hd0ef0284_0513eeff,
        64'hd0ef842a_e022e406,
        64'h1141d0cf_e06f6145,
        64'h64e26942_07848513,
        64'h864a6a02_69a270a2,
        64'h740285a2_d26fe0ef,
        64'h05048513_85ce8652,
        64'hd32fe0ef_85ca864e,
        64'h02848513_d3efe0ef,
        64'h05040993_02858913,
        64'h84aae44e_e84aec26,
        64'hf406842e_8652f022,
        64'h07858a13_e0527179,
        64'hd62fe06f_614564e2,
        64'h05048513_694269a2,
        64'h85ca864e_70a27402,
        64'hd7afe0ef_02840593,
        64'h864a0284_8513d88f,
        64'he0ef842e_05058913,
        64'h84aae84a_ec26f022,
        64'hf406864e_07858993,
        64'he44e7179_80826165,
        64'h7ae26a06_69a66946,
        64'h64e67406_70a6ffbf,
        64'hd0ef8556_002c8656,
        64'hd98ff0ef_8552002c,
        64'h865680ef_e0ef854a,
        64'h85d2864a_dacff0ef,
        64'h852685d2_864a822f,
        64'he0ef0028_85b20504,
        64'h0613decf_e0ef8556,
        64'h05098593_07840613,
        64'h07848a93_dfefe0ef,
        64'h854a85ca_864ee08f,
        64'he0ef8552_85a60289,
        64'h86130504_8a13deef,
        64'hf0ef854a_85d28622,
        64'h864fe0ef_84aa0285,
        64'h0913fc56_e8caeca6,
        64'hf4868622_89b285d2,
        64'he4ce0285_8a13842e,
        64'he0d2f0a2_71598082,
        64'h61657ae2_6a0669a6,
        64'h694664e6_740670a6,
        64'he30ff0ef_8556002c,
        64'h86568a6f_e0ef8552,
        64'h002c8656_8b0fe0ef,
        64'h854a85d2_864ae4ef,
        64'hf0ef8526_85d2864a,
        64'h8c4fe0ef_002885b2,
        64'h05040613_e8efe0ef,
        64'h85560509_85930784,
        64'h06130784_8a93ea0f,
        64'he0ef854a_85ca0289,
        64'h8613eacf_e0ef8552,
        64'h85a6864e_05048a13,
        64'he90ff0ef_854a85d2,
        64'h8622906f_e0ef84aa,
        64'h02850913_fc56e8ca,
        64'heca6f486_862289b2,
        64'h85d2e4ce_02858a13,
        64'h842ee0d2_f0a27159,
        64'hb7d5557d_bfe9d8df,
        64'he0ef8522_85a28082,
        64'h61116a4e_69ee790e,
        64'h74ae744e_70ee4501,
        64'hf0afe0ef_85a2864e,
        64'h07840513_02a78163,
        64'h839d01fa_4783a31f,
        64'hf0ef8522_f26fe0ef,
        64'h852285a2_02848613,
        64'he139a5df_f0ef1128,
        64'h97cfe0ef_010c0030,
        64'h1128c105_a6fff0ef,
        64'h1128f22f_f0ef010c,
        64'h00301128_f56fe0ef,
        64'h1810852e_010ce63f,
        64'he0ef0108_85a2f68f,
        64'he0ef8522_85a20030,
        64'hf72fe0ef_852285a2,
        64'h08b0ae0f_f0ef8522,
        64'h85a2f84f_e0ef8522,
        64'h85a20030_f8efe0ef,
        64'h852285a2_1810e9bf,
        64'he0ef8522_08acfa0f,
        64'he0ef852e_181008ac,
        64'headfe0ef_08a8180c,
        64'h9f4fe0ef_852e864a,
        64'h180cf92f_f0ef864a,
        64'h852e002c_fc6fe0ef,
        64'h1808002c_8626d624,
        64'h8493ed7f_e0ef0000,
        64'h14970028_85ce9f8f,
        64'he0ef854a_d8efe0ef,
        64'h8a2e0504_0913e9d2,
        64'hf1caf5a6_fd86854e,
        64'h842af9a2_02850993,
        64'hedce7111_80826165,
        64'h7ae26a06_69a66946,
        64'h64e67406_70a6feef,
        64'hf0ef8556_002c8656,
        64'ha64fe0ef_8552002c,
        64'h8656a6ef_e0ef854e,
        64'h85d2864e_80dff0ef,
        64'h852285d2_864ea82f,
        64'he0ef0028_85a28622,
        64'h84bfe0ef_85220504,
        64'h85930509_0613859f,
        64'he0ef8556_07890593,
        64'h07848613_07840a93,
        64'h86bfe0ef_854e85ce,
        64'h02890613_877fe0ef,
        64'h855285a2_864a0504,
        64'h0a1385bf_f0ef854e,
        64'h85d28626_ad0fe0ef,
        64'h02850993_842afc56,
        64'he4cef0a2_f4868626,
        64'h893285d2_e8ca0285,
        64'h8a1384ae_e0d2eca6,
        64'h71598082_61696baa,
        64'h6b4a6aea_7a0a79aa,
        64'h794a74ea_640e60ae,
        64'hbb8fe0ef_855208ac,
        64'h8656bc2f_e0ef855a,
        64'h180c8656_bccfe0ef,
        64'h854e002c_86562a81,
        64'hf87fe0ef_08a885d2,
        64'he58fe0ef_180885ce,
        64'he60fe0ef_002885da,
        64'hbf0fe0ef_855295a6,
        64'h864a3984_0593bfef,
        64'he0ef855a_95a6864a,
        64'h37040593_c0cfe0ef,
        64'h854e95a6_864a3484,
        64'h05930009_2913197d,
        64'hc20fe0ef_00894913,
        64'h855295a6_865e3204,
        64'h0593c32f_e0ef855a,
        64'h95a6865e_2f840593,
        64'hc40fe0ef_854e95a6,
        64'h865e2d04_0593000b,
        64'hab931bfd_c54fe0ef,
        64'h00794b93_855295a6,
        64'h865e2a84_0593c66f,
        64'he0ef855a_95a6865e,
        64'h28040593_c74fe0ef,
        64'h854e95a6_865e2584,
        64'h0593000b_ab931bfd,
        64'hc88fe0ef_00694b93,
        64'h855295a6_865e2304,
        64'h0593c9af_e0ef855a,
        64'h95a6865e_20840593,
        64'hca8fe0ef_854e95a6,
        64'h865e1e04_0593000b,
        64'hab931bfd_cbcfe0ef,
        64'h00594b93_855295a6,
        64'h865e1b84_0593ccef,
        64'he0ef855a_95a6865e,
        64'h19040593_cdcfe0ef,
        64'h854e95a6_865e1684,
        64'h0593000b_ab931bfd,
        64'hcf0fe0ef_00494b93,
        64'h855295a6_865e1404,
        64'h0593d02f_e0ef855a,
        64'h95a6865e_11840593,
        64'hd10fe0ef_854e95a6,
        64'h865e0f04_0593000b,
        64'hab931bfd_d24fe0ef,
        64'h00394b93_855295a6,
        64'h865e0c84_0593d36f,
        64'he0ef855a_95a6865e,
        64'h0a040593_d44fe0ef,
        64'h854e95a6_865e0784,
        64'h0593000b_ab931bfd,
        64'hd58fe0ef_00294b93,
        64'h855295a6_865e0504,
        64'h0593d6af_e0ef855a,
        64'h95a6865e_02840593,
        64'hd78fe0ef_854e865e,
        64'h009405b3_000bab93,
        64'hc88fe0ef_46648493,
        64'h041a0000_14971bfd,
        64'h8c058552_00449413,
        64'h00194b93_ccefe0ef,
        64'h05098a13_855a0ff9,
        64'h7913cdcf_e0ef03f6,
        64'h5a9384ae_02850b13,
        64'he55ee95a_ed5689aa,
        64'hf152f54e_fd26e1a2,
        64'h40f9093b_e5860017,
        64'h979b00f9_77b30ff6,
        64'h791343f6_5793f94a,
        64'h7155b7c1_00978023,
        64'hf96d0007_c503fcf8,
        64'h87e30785_00078023,
        64'ha03187b2_98be0016,
        64'h08939381_17824104,
        64'h07bbffe8_05e3fef6,
        64'h8fa3fe77_cce340f5,
        64'h07bbb775_0685fdc7,
        64'h1ce32705_00060023,
        64'hffd68fa3_01dfcb63,
        64'h00f50ebb_00e797bb,
        64'hfff68503_cf890006,
        64'h078302e3_04630605,
        64'h2805a029_40b2833b,
        64'h4705882e_8636ffe5,
        64'h89e38082_01416482,
        64'h6422ffe5_9be30685,
        64'heb812585_fff6c783,
        64'h0ff00413_53c51010,
        64'h02934e1d_4fbd4485,
        64'h10000f13_45810015,
        64'h0693fed7_91e30785,
        64'h00e60023_8b054107,
        64'h573b00f5_06330077,
        64'hf8130007_4703972e,
        64'h4037d71b_10000693,
        64'h4781e026_e4221141,
        64'h00003070_32635f30,
        64'h7032645f_30703266,
        64'h5f307032_615f3070,
        64'h326d5f30_70326934,
        64'h36767205_10040000,
        64'h002a0100_76637369,
        64'h72000000_34418082,
        64'h614500a0_35338d5d,
        64'h8d5970a2_8d5501f1,
        64'h47838d51_8d5d01e1,
        64'h470301d1_46838d59,
        64'h8d5501c1_460301b1,
        64'h47838d51_8d5d01a1,
        64'h47030191_46838d59,
        64'h8d550181_46030171,
        64'h47838d51_8d5d0161,
        64'h47030151_46838d59,
        64'h8d550141_46030131,
        64'h47838d51_8d5d0121,
        64'h47030111_46838d59,
        64'h8d550101_460300f1,
        64'h47838d51_8d5d00e1,
        64'h470300d1_46838d59,
        64'h8d5500c1_460300b1,
        64'h47838d51_8d5d00a1,
        64'h47030091_46838d59,
        64'h8d550081_46030071,
        64'h47838d51_8d5d0061,
        64'h47030051_46838d59,
        64'h8d550041_46030031,
        64'h47830021_47030001,
        64'h45030011_4683d53f,
        64'hf0eff406_850a85aa,
        64'h71798082_61458905,
        64'h70a20001_4503d6bf,
        64'hf0eff406_850a85aa,
        64'h71798082_61097d82,
        64'h7d227cc2_7c626b86,
        64'h6b266ac6_6a667986,
        64'h792674c6_01d50fa3,
        64'h00f50f23_00b50ea3,
        64'h01e50e23_00d50da3,
        64'h01050d23_01f50ca3,
        64'h00c50c23_01150ba3,
        64'h00e50b23_01c50823,
        64'h00550623_007504a3,
        64'h01550723_016506a3,
        64'h01750523_018503a3,
        64'h412ede9b_40c6d69b,
        64'h40d6561b_40aed79b,
        64'h402ed59b_012f6f33,
        64'h4046d81b_013fefb3,
        64'h4056589b_01476733,
        64'h00f50aa3_00b507a3,
        64'h010505a3_01150423,
        64'h4177571b_4146df1b,
        64'h41565f9b_4125d59b,
        64'h40b8581b_40d8d89b,
        64'h006e991b_47f200f5,
        64'h0a230046_999b0036,
        64'h1a1b47e2_00f509a3,
        64'h40a5da9b_4025db1b,
        64'h67c200f5_09234038,
        64'h5b9b4058_dc1b47b2,
        64'h00f508a3_74660085,
        64'h032347a2_006502a3,
        64'h40e3531b_01950223,
        64'h009501a3_01a50123,
        64'h01b500a3_00f50023,
        64'hce52cc7e_e87ac64e,
        64'hc44afc62_e0dee4da,
        64'h408e591b_410e599b,
        64'h0122e2b3_0133e3b3,
        64'h40775f9b_40f75a1b,
        64'h01efef33_01446433,
        64'h40635c9b_0154e4b3,
        64'h4087dd9b_4107dd1b,
        64'hf06ef46a_f8660017,
        64'h1f1b418e_5f9b4138,
        64'h529b4158_d39b4163,
        64'h541b4187_d49b0065,
        64'h991b0058_199b0038,
        64'h9a1b0023_1a9b01fe,
        64'hfeb30056_f6b301f6,
        64'h7633e8d6_ecd2f0ce,
        64'hf4ca01ee_8ebb01fe,
        64'h7e330057_77330055,
        64'hf5b301f8_78330058,
        64'hf8b301f3_73330057,
        64'hf7b341a6_de9b1ffd,
        64'h12fd0200_0fb70400,
        64'h02b79ea5_4196569b,
        64'h9e2141a7_561b0077,
        64'h073b419e_571b005e,
        64'h0e3b41a5_de1b01f5,
        64'h85bb4198_559b01d8,
        64'h083b41a8_d81b01c8,
        64'h88bb4193_589b0103,
        64'h033b41a7_d31b9fb1,
        64'h9f950027_979b9fb5,
        64'h0026979b_4196d69b,
        64'h01e686bb_41a6d69b,
        64'h9ea54196_d69b9ea1,
        64'h518441a6_d69bf8a6,
        64'h007686bb_4dc04196,
        64'hd69bfca2_005686bb,
        64'h711941a6_d69b0185,
        64'ha38301f6_86bb4196,
        64'hd69b0145_a28301d6,
        64'h86bb41a6_d69b0105,
        64'haf8301c6_86bb4196,
        64'hd69b00c5_ae830106,
        64'h86bb41a6_d69b0085,
        64'hae039eb1_4196d69b,
        64'h0045a803_9ebd41e6,
        64'h86bb0026_969b01e6,
        64'h86bb002f_169b0100,
        64'h07b74190_0245af03,
        64'h80826121_6b226ac2,
        64'h6a627982_792274c2,
        64'hd15cd118_cd540105,
        64'h2c2341f7_87bb4057,
        64'h073b4076_86bb7462,
        64'h4088083b_01152a23,
        64'h00652823_01c52623,
        64'h01d52423_c150c10c,
        64'h409888bb_41e585bb,
        64'h4123033b_413e0e3b,
        64'h415b063b_414e8ebb,
        64'h02462f83_02062283,
        64'h01c62383_4e00fc22,
        64'h4a44f826_418c0006,
        64'h2f0351dc_51984dd4,
        64'h0185a803_0145a883,
        64'h0105a303_00c5ae03,
        64'h0085ae83_00462a83,
        64'h01062903_00c62983,
        64'h0045ab03_00862a03,
        64'he45ae856_ec52f04e,
        64'hf44a7139_8082610d,
        64'h7ac664ca_c94cc91c,
        64'h01d52623_95c2407e,
        64'h8eb38f85_85e90153,
        64'hf3b38ced_95be97b2,
        64'h4193d793_93f69ebe,
        64'h078697c6_7b26646a,
        64'h97a20368_88b397fa,
        64'h02640433_692a97f2,
        64'h032f0f33_6d866cc6,
        64'h6c667a66_698ad158,
        64'hc15441f7_073303ca,
        64'h0e337622_c5104056,
        64'h06330092_f2b341a2,
        64'hde9300b6_02b39666,
        64'h06069676_025787b3,
        64'h96e286e9_015fffb3,
        64'h78420105_20234138,
        64'h08330096_f9b300b8,
        64'h06b39836_03b88eb3,
        64'h62a24058_0833080a,
        64'h98160022_9813419f,
        64'hd2930077_0fb3967e,
        64'h6d26976a_0706974e,
        64'h03640633_7b86410c,
        64'h0c330158_78334198,
        64'h5c93007c_08339c66,
        64'h0c069c42_037989b3,
        64'h977603b4_08339fb2,
        64'h02e88733_9e960373,
        64'h06339fb2_6bc203db,
        64'h8eb36de2_03b52023,
        64'h410d8db3_00987833,
        64'h41a85d13_00bd8833,
        64'h9dea0d86_9dc20327,
        64'h063392b2_03280833,
        64'h02c78633_78029c42,
        64'h03c282b3_76029fb2,
        64'h036f0c33_03478633,
        64'h986203cf_8fb39db2,
        64'h02670833_03ef0db3,
        64'h41b686b3_009dfdb3,
        64'h41addc93_00b68db3,
        64'h068696e6_9642033c,
        64'h8cb30287_08337ce2,
        64'h9c66032a_0cb396c2,
        64'h03f78c33_03bc8833,
        64'h96626de2_96ee03d8,
        64'h8c336cc2_01052e23,
        64'h41980833_015cfcb3,
        64'h419cdd13_00780cb3,
        64'h98660806_986a0367,
        64'h0db39662_03228d33,
        64'h02578633_986a038e,
        64'h0c3396b2_02ef0d33,
        64'h986a026e_863396b2,
        64'h03d98d33_032e0633,
        64'h983202d6_86b303c8,
        64'h8633cd10_03778833,
        64'h41a60633_009d7d33,
        64'h41ad5c93_00b60d33,
        64'h966e0606_9666966a,
        64'h02628cb3_9642032c,
        64'h0d33966a_02e80833,
        64'h03df0d33_966a6822,
        64'hf8424198_0833015c,
        64'hfcb3419c_dd930078,
        64'h0cb39866_0806986e,
        64'h028e0d33_026c0db3,
        64'h986a0317_8633986e,
        64'h03288d33_f43241a6,
        64'h0633009d_7d3341ad,
        64'h5c9300b6_0d3303dd,
        64'h0db30606_96666d22,
        64'h986a036b_8cb30337,
        64'h8833fc66_03cf0d33,
        64'h033c8cbb_966a037c,
        64'h8b3b966e_02680d33,
        64'hfe000ab7_966a0324,
        64'h0db3f8d6_010003b7,
        64'h001b9c1b_ece2fc00,
        64'h04b7e826_020005b7,
        64'hec2e966e_034a0d33,
        64'h001f149b_001a1e9b,
        64'he9264115_85bb0025,
        64'h959b0115_85bb0028,
        64'h959bf4da_0018981b,
        64'h03e78633_4053033b,
        64'h0023131b_01c5ab83,
        64'h0019941b_f0deed22,
        64'h0053033b_0022931b,
        64'h0185a883_02ee0db3,
        64'h0145a983_e14e0205,
        64'ha283e4ea_e0ee0016,
        64'h979b0017_171bf03e,
        64'he43a02fc_893b001f,
        64'h9e1be54a_02600c93,
        64'h0085aa03_e8e6fcd2,
        64'h0105af03_71354194,
        64'h45d80045_af8351dc,
        64'h8082610d_690a64aa,
        64'h644a60ea_b56ff0ef,
        64'h854a002c_8626a63f,
        64'hf0ef852e_002ca6bf,
        64'hf0ef852e_002cb70f,
        64'hf0ef180c_85320030,
        64'hf87da7ff_f0ef852e,
        64'h347d180c_03100413,
        64'ha8dff0ef_852e180c,
        64'hb92ff0ef_08ac8532,
        64'h1810f87d_aa1ff0ef,
        64'h852e347d_08ac0630,
        64'h0413aaff_f0ef08a8,
        64'h180cbb4f_f0ef0030,
        64'h852e180c_f87dac3f,
        64'hf0ef852e_347d180c,
        64'h03100413_ad1ff0ef,
        64'h1808002c_bd6ff0ef,
        64'h180c8532_0030f87d,
        64'hae5ff0ef_852e347d,
        64'h180c4425_af1ff0ef,
        64'h852e180c_bf6ff0ef,
        64'h08ac8532_1810f87d,
        64'hb05ff0ef_852e347d,
        64'h08ac444d_b11ff0ef,
        64'h08a8180c_c16ff0ef,
        64'h0030852e_180cf87d,
        64'hb25ff0ef_852e347d,
        64'h180c4425_b31ff0ef,
        64'h1808002c_c36ff0ef,
        64'h180c8532_0030f87d,
        64'hb45ff0ef_852e347d,
        64'h180c4411_b51ff0ef,
        64'h1808002c_c56ff0ef,
        64'h180c8532_0030b63f,
        64'hf0ef852e_002cc68f,
        64'hf0ef852e_1810002c,
        64'hc72ff0ef_85a68532,
        64'h1810b7ff_f0ef852e,
        64'h180cb87f_f0ef1808,
        64'h002cb8ff_f0ef84ae,
        64'he526e922_ed060028,
        64'h892ae14a_71358082,
        64'h612974aa_744a70ea,
        64'hcaaff0ef_8526102c,
        64'h860af87d_bb9ff0ef,
        64'h852e347d_102c4411,
        64'hbc5ff0ef_852e102c,
        64'hccaff0ef_088c8532,
        64'h1030f87d_bd9ff0ef,
        64'h852e347d_088c0310,
        64'h0413be7f_f0ef852e,
        64'h088ccecf_f0ef18ac,
        64'h85320890_f87dbfbf,
        64'hf0ef852e_347d18ac,
        64'h06300413_c09ff0ef,
        64'h18a8088c_d0eff0ef,
        64'h1030852e_088cf87d,
        64'hc1dff0ef_852e347d,
        64'h088c0310_0413c2bf,
        64'hf0ef0888_102cd30f,
        64'hf0ef088c_85321030,
        64'hf87dc3ff_f0ef852e,
        64'h347d088c_4425c4bf,
        64'hf0ef852e_088cd50f,
        64'hf0ef18ac_85320890,
        64'hf87dc5ff_f0ef852e,
        64'h347d18ac_444dc6bf,
        64'hf0ef18a8_088cd70f,
        64'hf0ef1030_852e088c,
        64'hf87dc7ff_f0ef852e,
        64'h347d088c_4425c8bf,
        64'hf0ef0888_102cd90f,
        64'hf0ef088c_85321030,
        64'hf87dc9ff_f0ef852e,
        64'h347d088c_4411cabf,
        64'hf0ef0888_102cdb0f,
        64'hf0ef0890_852e102c,
        64'hcbdff0ef_0888858a,
        64'hdc2ff0ef_850a858a,
        64'h1030dccf_f0ef8532,
        64'h85a21030_cd9ff0ef,
        64'h852e102c_ce1ff0ef,
        64'h1028858a_ce9ff0ef,
        64'h842ef922_fd06850a,
        64'h84aaf526_71318082,
        64'h610d7ac6_64cac94c,
        64'hc91c01c5_262395f6,
        64'h407e0e33_8f8585e9,
        64'h0153f3b3_8ced95be,
        64'h97b24193_d79393f2,
        64'h9e3e97c2_7b26646a,
        64'h97a20368_083397fa,
        64'h03140433_6d26692a,
        64'h979a032f_0f336c66,
        64'h7a66698a_01f52223,
        64'hc1149fea_413686b3,
        64'h41afdf93_009ff9b3,
        64'h026a0333_00b68fb3,
        64'h7622c510_40560633,
        64'h0092f2b3_41a2de13,
        64'h00b602b3_96629672,
        64'h03f787b3_6d8603b8,
        64'h0e336fa2_96fe405f,
        64'h8fb30f8a_9f960022,
        64'h9f93967e_6cc6d158,
        64'h7ec241d7_0733015e,
        64'hfeb3419e_d2930077,
        64'h0eb39766_974e0364,
        64'h06337b86_97720379,
        64'h89b341dd_0d33015e,
        64'hfeb3419e_dc13007d,
        64'h0eb39d62_9d7602e8,
        64'h07339fb2_03b40eb3,
        64'h9e160378_86339fb2,
        64'h6bc203cb_8e336de2,
        64'h03b52023_41dd8db3,
        64'h009efeb3_41aedc93,
        64'h00bd8eb3_9de69df6,
        64'h03270633_92b2032e,
        64'h8eb302c7_86337e82,
        64'h9d760262_82b37602,
        64'h9fb2036f_0d330347,
        64'h86339eea_026f8fb3,
        64'h9db20317_0eb303ef,
        64'h0db341b6_86b3009d,
        64'hfdb341ad_dc1300b6,
        64'h8db396e2_9676033c,
        64'h0c330287_0eb37c62,
        64'h9d6203f7_8d3396f6,
        64'h032a0c33_03bd0eb3,
        64'h96626de2_96ee03c8,
        64'h0c336d42_01d52e23,
        64'h41ae8eb3_015d7d33,
        64'h419d5c93_007e8d33,
        64'h9ee69eea_03670db3,
        64'h96620322_8d330257,
        64'h86339eea_03830c33,
        64'h96b202ef_0d339eea,
        64'h031e0633_96b203c9,
        64'h8d330323_06339eb2,
        64'h02d686b3_02680633,
        64'hcd100377_8eb341a6,
        64'h0633009d_7d3341ad,
        64'h5c9300b6_0d33966e,
        64'h9666966a_03128cb3,
        64'h9676032c_0d3302ee,
        64'h8eb3966a_6ea2f876,
        64'h419e8eb3_015cfcb3,
        64'h419cdd93_007e8cb3,
        64'h9ee69eee_03cf0d33,
        64'h966a031c_0db30283,
        64'h0d339eea_03078633,
        64'h9eee0328_0d33f432,
        64'h41a60633_009d7d33,
        64'h41ad5c93_00b60d33,
        64'h03cd0db3_96666d22,
        64'h9eea036b_8cb30337,
        64'h8eb3fc66_026f0d33,
        64'h033c8cbb_966a037c,
        64'h8b3b966e_031e8d33,
        64'hfe000ab7_966a0324,
        64'h0db3f8d6_010003b7,
        64'h001b9c1b_ece2fc00,
        64'h04b7e826_020005b7,
        64'hec2e966e_034a0d33,
        64'h001f149b_001a1e1b,
        64'he9264105_85bb0025,
        64'h959b0105_85bb0028,
        64'h159bf4da_00181e9b,
        64'h03e78633_01c5ab83,
        64'h405888bb_f0de0019,
        64'h941b0028_989bed22,
        64'h005888bb_0022989b,
        64'h0185a803_02e30db3,
        64'h0145a983_e14e0205,
        64'ha283e4ea_e0ee0016,
        64'h979b0017_171bf03e,
        64'he43a02fc_893b001f,
        64'h931be54a_02600c93,
        64'h0085aa03_e8e6fcd2,
        64'h0105af03_71354194,
        64'h45d80045_af8351dc,
        64'h8082d15c_d118cd54,
        64'hcd100105_2a230115,
        64'h28230065_262301c5,
        64'h242301d5_2223c10c,
        64'h40b005bb_40f007bb,
        64'h40e0073b_40d006bb,
        64'h40c0063b_4100083b,
        64'h411008bb_4060033b,
        64'h41c00e3b_41d00ebb,
        64'h418c51dc_51984dd4,
        64'h4d900145_a8030105,
        64'ha88300c5_a3030085,
        64'hae030045_ae838082,
        64'h61456a82_6a22d15c,
        64'hd11897ae_8f1187e9,
        64'h8e7d97ba_01fe8733,
        64'h69c2cd54_01052c23,
        64'h96fa86e9_40e80833,
        64'h00c6f733_00f806b3,
        64'h981e02ef_8fb36962,
        64'h01152823_406888b3,
        64'hc9549696_86e900c6,
        64'hf33300f8_86b398ca,
        64'h02e383b3_74820065,
        64'h2423c554_41c30333,
        64'h96a686e9_00c6fe33,
        64'h00f306b3_935202e9,
        64'h09337422_01c52023,
        64'hc154408e_0e3396ce,
        64'h86e900c6_f43300fe,
        64'h06b39e56_02ea0a33,
        64'h40df0f33_8ee14196,
        64'hde9396fa_02ea8ab3,
        64'h41d282b3_008efeb3,
        64'h419ed813_00d28eb3,
        64'h02ef0f33_fc000637,
        64'h410484b3_00887833,
        64'h41985893_00d48833,
        64'h02e282b3_020007b7,
        64'h40fe0e33_411e85b3,
        64'h0e0a0205_af834109,
        64'h89b30088_78334198,
        64'h531300d9_883302e4,
        64'h84b39e3e_0088f8b3,
        64'h00279e13_0185a383,
        64'hfe000437_4198d793,
        64'hf42200de_88b30105,
        64'ha90302e9_89b30100,
        64'h06b7ec4a_0085aa03,
        64'he4520005_aa83e056,
        64'h01c5af03_0145a283,
        64'h45c402ee_8eb3f026,
        64'hb4270713_0045a983,
        64'h6779e84e_0245ae83,
        64'h71798082_61516bce,
        64'h7a8e79ce_796ec94c,
        64'hc918c554_8e9d95de,
        64'h41270733_85e90137,
        64'hf7b30125_f93395ba,
        64'h97564197_d7130076,
        64'h87b300f8_06b397b6,
        64'h6bea6aca_97ba035b,
        64'h86b36b6e_643297fa,
        64'h028b0733_7dca7d6a,
        64'h6c8e6c2e_7a2e6492,
        64'h97f6034c_8f33c510,
        64'h41c60633_012e7e33,
        64'hd1580115_22239896,
        64'hc11441a8_d89341f6,
        64'h86b303dd_0eb30128,
        64'hffb397fe_41ae5813,
        64'h00b60e33_40670733,
        64'h01337333_fe0009b7,
        64'h964e00b6_88b39646,
        64'h96c203b7_87b341c8,
        64'h0833080a_9872002e,
        64'h18134193_5e130077,
        64'h03330100_03b7971e,
        64'h977a0308_88b378a6,
        64'h9646035f_0f336862,
        64'h9742028b_8633989a,
        64'h02880833_6d229772,
        64'h03ab08b3_9fb2034e,
        64'h0e339fc6_02960633,
        64'h7b86935e_038f0fb3,
        64'h67827b22_405f82b3,
        64'h00f2f2b3_4192d993,
        64'h92fe03dc_83330100,
        64'h02b79fda_9f96fe00,
        64'h07b7971a_035782b3,
        64'h03d70733_7ae698d6,
        64'h03352023_6ce64059,
        64'h89b30122_f2b341a2,
        64'hd39300b9_82b399e6,
        64'h99960318_08b30276,
        64'h02b39f96_63e29b9e,
        64'h028f8fb3_6a267fa6,
        64'h027a03b3_9afe63c2,
        64'h931e02ef_8fb36a22,
        64'h99d203b3_83b3028f,
        64'h09b36d86_03be0ab3,
        64'h9bd692ce_029b8bb3,
        64'h6b8240db_86b30126,
        64'hf6b341a6_db13025b,
        64'h02b300bb_86b39bb6,
        64'h62a67b06_931602db,
        64'h06b30293_03337b0a,
        64'h9a5a7dc6_9b6e03a8,
        64'h0a3366e2_9ab603de,
        64'h0b3399d2_7d4203a6,
        64'h0ab396da_03d989b3,
        64'h9bd6031f_06b379a2,
        64'h92ce02f4_0bb30389,
        64'h89b30175_2e23678a,
        64'h7c62418b_8bb300fc,
        64'h7c33419c_5c93fe00,
        64'h07b79c5e_01000c37,
        64'h9bbe9be2_77aa0397,
        64'h8c339a62_9ab67ce6,
        64'h034c8a33_67826a06,
        64'h6ce602fc_8ab392d2,
        64'h7cc29de6_031282b3,
        64'h9bd603b7_0db30286,
        64'h0bb36dc2_9b6e03cf,
        64'h8b330378_0db396da,
        64'h7b829c5e_02de86b3,
        64'h7686029c_0c339cb6,
        64'h6c229a62_02938cb3,
        64'h77a603f7_8c3303ba,
        64'h0a339ae2_9be6035f,
        64'h0ab367aa_03778bb3,
        64'h6aa69b56_7dc696ee,
        64'h7be2037b_0b336782,
        64'h03a306b3_7ba29c5e,
        64'hf53ecd14_6b424166,
        64'h86b3012b_7b3341ab,
        64'h579300b6_8b3396be,
        64'h96da03d8_0c336d46,
        64'h9ce2036d_0b336b62,
        64'h9ada0316_0cb36d22,
        64'h9de603a4_8ab39bd6,
        64'h03198db3_96ee037e,
        64'h0bb36d66_6b869c5e,
        64'h028d0db3_03bf0bb3,
        64'h9b5e030f_8c336d02,
        64'h9ce2037d_0bb3034f,
        64'h8cb36ba2_03728c33,
        64'h96e296e6_03860c33,
        64'h7b829ade_03df0cb3,
        64'h7c420297_0bb39ae2,
        64'h9b5e0383_8c336d46,
        64'h9b6603a8_8bb303ef,
        64'h8b3396da_6d0202cd,
        64'h0cb37dc6_ed5e9ae6,
        64'h03680b33_7c62418b,
        64'h8bb301bc_7c33419c,
        64'h5793fe00_0db79c5e,
        64'h01000c37_9be29bee,
        64'h03130cb3_9be603b7,
        64'h8db3ecbe_7de67d02,
        64'h6b429ada_028c8cb3,
        64'h03b98b33_6ca29be6,
        64'h025f8ab3_96da039d,
        64'h0cb3e956_029e0b33,
        64'h416a8ab3_012b7b33,
        64'h41ab5c13_96e26d02,
        64'h00ba8b33_9ada03a7,
        64'h0c336ca6_9ae2036c,
        64'h8b336d46_6b629bda,
        64'h028d0c33_9be203d6,
        64'h0b337ca2_96da039f,
        64'h0c3396e2_03138b33,
        64'h9ada033f_86b36c86,
        64'h036c8b33_9ab67b42,
        64'h03630c33_87ea03d7,
        64'h86b39ab6_7b029bda,
        64'h02d606b3_02980b33,
        64'h9bda66c2_9ab6038e,
        64'h0b33fc00_09376ca2,
        64'he16641c9_0cbb0029,
        64'h191b9bda_029f0ab3,
        64'h01c9093b_002e191b,
        64'h96caf4d6_40ea8abb,
        64'h002a9a9b_00ea8abb,
        64'h00271a9b_96d60317,
        64'h0b33f8ee_020005b7,
        64'hf12e4105_85bb0025,
        64'h959b0105_85bb0028,
        64'h159b9bda_031e0ab3,
        64'h8de6fcee_6782f0be,
        64'h407587bb_e03e0025,
        64'h959b4147_87bb0027,
        64'h979b026f_8bb30075,
        64'h85bb0023_959b0147,
        64'h87bbec2e_002a179b,
        64'h7c62e462_405c0c3b,
        64'h002c1c1b_03938b33,
        64'h005c0c3b_00229c1b,
        64'he856000b_859b96da,
        64'hf42e001d_9b9b413b,
        64'h8d3b4065_85bb03a8,
        64'h0933e8ea_f84a0025,
        64'h959b0019_191b002b,
        64'h9b9be4ca_001c1d1b,
        64'h006585bb_013b8bbb,
        64'h0023159b_51800029,
        64'h9b9b0004_0a9be55e,
        64'h8dd64176_063b0026,
        64'h161b001d_941b0176,
        64'h063b0245_aa83e0ee,
        64'h002b961b_01c5a903,
        64'h02062a03_01c62283,
        64'h01862983_01462303,
        64'h0185ae83_00062f03,
        64'h0085a883_49840086,
        64'h2e030046_2803027f,
        64'h86b3f022_fc62fd6a,
        64'hf1d6f5d2_f9cefdca,
        64'he2260145_ad830287,
        64'h0b330246_2b83f96e,
        64'he9deedda_00c5ac03,
        64'h001c941b_e5e2e622,
        64'h01062383_0005af83,
        64'h46580045_ac83e1e6,
        64'h716d8082_610d6d86,
        64'h6d266cc6_6c667b86,
        64'h7b267ac6_7a66698a,
        64'h692a64ca_d15cd10c,
        64'hcd140145_2a2397f6,
        64'h40bf05b3_411986b3,
        64'h9a1687e9_41aa5a13,
        64'h646a4053_82b3cd40,
        64'h8dfdc910_01052423,
        64'h01f52023_40c30633,
        64'h01652623_01752223,
        64'h943a97fa_410e0833,
        64'h846900ba_763340da,
        64'h8fb340e6_073301f2,
        64'hf2b39b26_9bca00b4,
        64'h78b341ab_db9300bb,
        64'hf6b341ab_5b1341d6,
        64'h8eb300bb_783301f7,
        64'h77334098_04b34128,
        64'h893300f3_0a3300f9,
        64'h843301f4_f4b301f9,
        64'h793300fe_0b3301fe,
        64'hfeb3935a_fc0005b7,
        64'h00fa8bb3_01a58f33,
        64'h99d24192_d9934194,
        64'hd3130d12_0a1e9e5e,
        64'h41975593_00231b13,
        64'h9afafe00_0fb74199,
        64'h5e13408a_8ab300bd,
        64'h6d33016a_6a33005e,
        64'h1b9301bf_6f339732,
        64'h01736333_00e382b3,
        64'h00e804b3_0a8a0f62,
        64'h01aced33_0149ea33,
        64'h0064e333_018e6e33,
        64'h01fdedb3_0616080e,
        64'h00e88933_0dc20d42,
        64'h0a420342_9aa201c9,
        64'h6e330ca2_09a204a2,
        64'h005fefb3_089a0e42,
        64'h00241a93_0fa20156,
        64'h663301a5_c5830922,
        64'h0145cb03_00d5cb83,
        64'h419ed413_0035cf03,
        64'h0075cc03_79c262e2,
        64'h01386833_0053e3b3,
        64'h7a6200e6_8eb30025,
        64'hcd8301c5_cd0301b5,
        64'hcc8300f5_c30303e2,
        64'hec76fc5e_f85a6a82,
        64'h01000737_e06269a2,
        64'h0138e8b3_0158e8b3,
        64'h73a20005_ce830072,
        64'he2b301d6_f6b30165,
        64'hcb830155_cb0302c2,
        64'h08a2068a_0ac20143,
        64'he3b3ffc7_8e93f47a,
        64'h0175cc03_69c203a2,
        64'h00c9e633_020007b7,
        64'h064209a2_7a020135,
        64'hcf0300e5_c4830148,
        64'h6833e426_e822f03a,
        64'h0095ce03_0085c903,
        64'h0015cf83_0125c283,
        64'h0065ca83_0055c883,
        64'h08220a42_0115c383,
        64'h0195c603_0185c983,
        64'h0105c703_8ed900a5,
        64'hc4830045_c4038edd,
        64'h00c5ca03_00b5c803,
        64'h07a206c2_01d5c703,
        64'h01e5c783_01f5c683,
        64'hf8d6fcd2_e14ee54a,
        64'he926ed22_e0eee4ea,
        64'he8e6ece2_f0def4da,
        64'h71358082_d15cd118,
        64'hcd54cd10_01052a23,
        64'h01152823_00652623,
        64'h01c52423_01d52223,
        64'h01e52023_51dc5198,
        64'h4dd44d90_0145a803,
        64'h0105a883_00c5a303,
        64'h0085ae03_0045ae83,
        64'h0005af03_80826149,
        64'h7dc27d62_6c866c26,
        64'h6bc66b66_7a867a26,
        64'h79c67966_648ad1d4,
        64'hd1900104_c633642a,
        64'h8ea1cdc8_0065ac23,
        64'h01c5aa23_01d5a823,
        64'hc5dcc598_0055a223,
        64'h0075a023_01e7c7b3,
        64'h01f74733_00664333,
        64'h01b3c3b3_64a26442,
        64'h01144533_d1440325,
        64'h20230135_2e230145,
        64'h2c230155_2a230165,
        64'h28230175_26230185,
        64'h24230195_222301a5,
        64'h20230109_49330119,
        64'hc9b301eb_cbb301fc,
        64'h4c338cb5_006a4a33,
        64'h01bd4d33_762201c6,
        64'h4e3301ca_cab36402,
        64'h0082c2b3_760201d6,
        64'h4eb3008c_ccb301db,
        64'h4b336662_8ef10106,
        64'h78330116_78b30066,
        64'h733301c6_7e3301d6,
        64'h7eb301e6_7f3301f6,
        64'h7fb38c71_01b67db3,
        64'h8ea50109_483300fb,
        64'hcf3300ec_4fb3005c,
        64'hc433007d_4db340c0,
        64'h063b66c2_00d9c8b3,
        64'h6822011a_4333010a,
        64'hce33f446_f0425144,
        64'h02052903_6682ec36,
        64'h01c52983_00db4eb3,
        64'he81ae426_e02245dc,
        64'h45980045_a2830005,
        64'ha3830185_2a030145,
        64'h2a8300c5_2b830085,
        64'h2c030045_2c830005,
        64'h2d030185_a8830145,
        64'ha803f8ce_f86efc6a,
        64'he0e6e4e2_e8def0d6,
        64'hf4d2fcca_0245a303,
        64'h51844dc0_01052b03,
        64'h4994ecda_e126e522,
        64'h71758082_61216b82,
        64'h6b226ac2_6a627982,
        64'h792274c2_03e52223,
        64'h03f52023_00552e23,
        64'h00752c23_00ff4f33,
        64'h00efcfb3_00d2c2b3,
        64'h00b3c3b3_7462c940,
        64'hc904c110_01252623,
        64'h01352423_01452223,
        64'h01044433_0114c4b3,
        64'h00694933_01c9c9b3,
        64'h01da4a33_00cb4633,
        64'h01567633_8ff18f71,
        64'h8ef18df1_01067833,
        64'h011678b3_00667333,
        64'h01c67e33_01d67eb3,
        64'h00ff47b3_00efc733,
        64'h00d2c6b3_01044833,
        64'h0114c8b3_00694333,
        64'h01c9ce33_01da4eb3,
        64'h015b4ab3_0173c5b3,
        64'h40c0063b_02452f03,
        64'h02052f83_01c52283,
        64'h01852383_49404904,
        64'h00c52903_00852983,
        64'h00452a03_00052b03,
        64'h0005aa83_51dc5198,
        64'h4dd40185_ab830145,
        64'ha8030105_a88300c5,
        64'ha3030085_ae030045,
        64'hae83e05e_e45ae856,
        64'hec52f04e_f44af826,
        64'hfc227139_80826121,
        64'h6b226ac2_6a627982,
        64'h792274c2_d15cd118,
        64'hcd540105_2c2301f7,
        64'h87bb0057_073b0076,
        64'h86bb7462_0088083b,
        64'h01152a23_00652823,
        64'h01c52623_01d52423,
        64'hc150c10c_009888bb,
        64'h01e585bb_0123033b,
        64'h013e0e3b_015b063b,
        64'h014e8ebb_525c5218,
        64'h4e540186_28030146,
        64'h2883420c_0005af03,
        64'h0245af83_0205a283,
        64'h01c5a383_01062303,
        64'h00c62e03_00862e83,
        64'h00462b03_4d8049c4,
        64'h0105a903_00c5a983,
        64'h0085aa03_0045aa83,
        64'he45ae856_ec52f04e,
        64'hf44af826_fc227139,
        64'h80820205_22230205,
        64'h20230005_2e230005,
        64'h2c230005_2a230005,
        64'h28230005_26230005,
        64'h24230005_2223c11c,
        64'h47858082_02052223,
        64'h02052023_00052e23,
        64'h00052c23_00052a23,
        64'h00052823_00052623,
        64'h00052423_00052223,
        64'h00052023_00003070,
        64'h32635f30_7032645f,
        64'h30703266_5f307032,
        64'h615f3070_326d5f30,
        64'h70326934_36767205,
        64'h10040000_002a0100,
        64'h76637369_72000000,
        64'h3441b7c5_fcc89ee3,
        64'h080500f8_00230505,
        64'h08850008_c7838082,
        64'h40010113_fcaefce3,
        64'h400e0e13_00678963,
        64'h00084783_fec718e3,
        64'h0785fed7_0fa300b7,
        64'h80230705_0007c683,
        64'h87f2870a_888a8872,
        64'hfffece93_0aa00313,
        64'hfaa00593_45014001,
        64'h06138e2a_80000eb7,
        64'hc0010113_00003070,
        64'h32635f30_7032645f,
        64'h30703266_5f307032,
        64'h615f3070_326d5f30,
        64'h70326934_36767205,
        64'h10040000_002a0100,
        64'h76637369_72000000,
        64'h34418082_00f68023,
        64'h0ff7f793_8fd900a7,
        64'h173b4705_0006c783,
        64'h400006b7_808200e6,
        64'h80238f7d_fff7c793,
        64'h00a797bb_47850006,
        64'hc7034000_06b78082,
        64'h00e78623_477d0007,
        64'h82234000_07b78082,
        64'h00054503_808200b5,
        64'h00230030_7032635f,
        64'h30703264_5f307032,
        64'h665f3070_32615f30,
        64'h70326d5f_30703269,
        64'h34367672_05100400,
        64'h00002a01_00766373,
        64'h69720000_00344100,
        64'h0a0d2165_6e6f6420,
        64'h00000020_6567616d,
        64'h6920746f_6f622067,
        64'h6e697970_6f630a0d,
        64'h00000000_2d2d2d2d,
        64'h2d2d2d2d_2d2d2d2d,
        64'h2d2d2d2d_2d2d2d2d,
        64'h2d2d2d2d_2d2d0a0d,
        64'h0000203a_657a6569,
        64'h735f6174_61640a0d,
        64'h00000000_00000020,
        64'h3a61626c_5f747361,
        64'h6c5f6174_61640a0d,
        64'h00000000_0000203a,
        64'h61626c5f_74737269,
        64'h665f6174_61640a0d,
        64'h00000000_00000009,
        64'h3a656d61_6e090a0d,
        64'h00093a73_65747562,
        64'h69727474_61090a0d,
        64'h00000009_3a61626c,
        64'h20747361_6c090a0d,
        64'h0000093a_61626c20,
        64'h74737269_66090a0d,
        64'h00000000_00000000,
        64'h09202020_20203a64,
        64'h69756720_6e6f6974,
        64'h69747261_70090a0d,
        64'h00000000_00000000,
        64'h093a6469_75672065,
        64'h70797420_6e6f6974,
        64'h69747261_70090a0d,
        64'h00000000_20797274,
        64'h6e65206e_6f697469,
        64'h74726170_20747067,
        64'h00000009_20203a73,
        64'h65697274_6e65206e,
        64'h6f697469_74726170,
        64'h20657a69_73090a0d,
        64'h00000009_3a736569,
        64'h72746e65_206e6f69,
        64'h74697472_61702072,
        64'h65626d75_6e090a0d,
        64'h00000009_2020203a,
        64'h61626c20_73656972,
        64'h746e6520_6e6f6974,
        64'h69747261_70090a0d,
        64'h00093a61_646c2070,
        64'h756b6361_62090a0d,
        64'h00000000_00000000,
        64'h093a6162_6c20746e,
        64'h65727275_63090a0d,
        64'h00000009_3a646576,
        64'h72657365_72090a0d,
        64'h00093a72_65646165,
        64'h685f6372_63090a0d,
        64'h00000000_00000909,
        64'h3a657a69_73090a0d,
        64'h00000009_3a6e6f69,
        64'h73697665_72090a0d,
        64'h0000093a_65727574,
        64'h616e6769_73090a0d,
        64'h00000000_003a7265,
        64'h64616568_20656c62,
        64'h6174206e_6f697469,
        64'h74726170_20747067,
        64'h0000203a_65756c61,
        64'h76206e72_75746572,
        64'h2079706f_63206473,
        64'h00000000_0000000a,
        64'h0d216465_6c696166,
        64'h20647261_63204453,
        64'h00000000_0000000a,
        64'h0d216465_7a696c61,
        64'h6974696e_69206473,
        64'h00000000_0a0d676e,
        64'h69746978_65202e2e,
        64'h2e647320_657a696c,
        64'h61697469_6e692074,
        64'h6f6e2064_6c756f63,
        64'hb7a954f9_b58ff0ef,
        64'h6a050513_fffff517,
        64'hbf6ff0ef_8526b6af,
        64'hf0ef07a5_05130000,
        64'h0517b76f_f0ef06e5,
        64'h05130000_0517bfa5,
        64'h54f9b86f_f0ef6ce5,
        64'h0513ffff_f517c24f,
        64'hf0ef8556_b98ff0ef,
        64'h0a850513_00000517,
        64'hba4ff0ef_09c50513,
        64'h00000517_b75d54f9,
        64'hbb4ff0ef_6fc50513,
        64'hfffff517_c52ff0ef,
        64'h8526bc6f_f0ef0d65,
        64'h05130000_0517bd2f,
        64'hf0ef0ca5_05130000,
        64'h0517bfd1_54fdbe2f,
        64'hf0ef09a5_05130000,
        64'h05178082_61616c02,
        64'h6ba26b42_6ae27a02,
        64'h79a27942_74e26406,
        64'h852660a6_fb040113,
        64'hc0cff0ef_33c50513,
        64'h00000517_ed1584aa,
        64'hba7ff0ef_9e0d2605,
        64'h8562020b_2583028b,
        64'h3603c2ef_f0ef3465,
        64'h05130000_0517c3af,
        64'hf0ef3325_05130000,
        64'h0517cd8f_f0ef40a7,
        64'h85330785_020b3503,
        64'h028b3783_c58ff0ef,
        64'h34050513_00000517,
        64'hcf6ff0ef_028b3503,
        64'hc6cff0ef_33c50513,
        64'h00000517_d0aff0ef,
        64'h020b3503_c80ff0ef,
        64'h33850513_00000517,
        64'hf37a9fe3_080a0a13,
        64'h08098993_08048913,
        64'hc9cff0ef_2a857e65,
        64'h0513ffff_f517ff24,
        64'h9be3d8ef_f0ef0485,
        64'h0004c503_cb8ff0ef,
        64'h36050513_00000517,
        64'hd56ff0ef_0109b503,
        64'hcccff0ef_36450513,
        64'h00000517_d6aff0ef,
        64'h0089b503_ce0ff0ef,
        64'h36850513_00000517,
        64'hd7eff0ef_fb890493,
        64'h0009b503_cf8ff0ef,
        64'h37050513_00000517,
        64'hff349be3_de8ff0ef,
        64'h04850004_c50384d2,
        64'hd14ff0ef_36c50513,
        64'h00000517_ff449be3,
        64'he04ff0ef_04850004,
        64'hc503f809_0493d32f,
        64'hf0ef36a5_05130000,
        64'h0517e1ef_f0ef0ffa,
        64'hf513d46f_f0ef3665,
        64'h05130000_05174b91,
        64'h01010a13_02010993,
        64'h08010913_1a051a63,
        64'h8aaa8b0a_cf3ff0ef,
        64'h850a4605_71010489,
        64'h2583d76f_f0ef8be5,
        64'h05130000_0517dc8f,
        64'hf0ef4556_d88ff0ef,
        64'h38850513_00000517,
        64'hddaff0ef_4546d9af,
        64'hf0ef37a5_05130000,
        64'h0517e38f_f0ef6526,
        64'hdacff0ef_36c50513,
        64'h00000517_e4aff0ef,
        64'h7502dbef_f0ef36e5,
        64'h05130000_0517e5cf,
        64'hf0ef6562_dd0ff0ef,
        64'h36850513_00000517,
        64'he22ff0ef_4552de2f,
        64'hf0ef36a5_05130000,
        64'h0517e34f_f0ef4542,
        64'hdf4ff0ef_36c50513,
        64'h00000517_e46ff0ef,
        64'h4532e06f_f0ef36e5,
        64'h05130000_0517e58f,
        64'hf0ef4522_e18ff0ef,
        64'h37050513_00000517,
        64'heb6ff0ef_6502e2af,
        64'hf0ef3725_05130000,
        64'h0517e36f_f0ef35e5,
        64'h05130000_05172c05,
        64'h126384aa_890add5f,
        64'hf0ef850a_45854605,
        64'h7101e56f_f0ef3365,
        64'h05130000_05172605,
        64'h1c63ce1f_f0ef8c2a,
        64'h0880e45e_e85aec56,
        64'hf052f44e_f84afc26,
        64'he486e062_e0a2715d,
        64'h00003070_32635f30,
        64'h7032645f_30703266,
        64'h5f307032_615f3070,
        64'h326d5f30_70326934,
        64'h36767205_10040000,
        64'h002a0100_76637369,
        64'h72000000_3441002e,
        64'h00000000_0000000a,
        64'h0d6b636f_6c622044,
        64'h53206461_65722074,
        64'h6f6e2064_6c756f63,
        64'h0000000a_0d202e2e,
        64'h2e445320_676e697a,
        64'h696c6169_74696e69,
        64'h00000031_34646d63,
        64'h00000035_35646d63,
        64'h00000000_30646d63,
        64'h00000020_3a206573,
        64'h6e6f7073_65720920,
        64'h00000000_0020646e,
        64'h616d6d6f_63204453,
        64'h00000000_0000b7f1,
        64'h547df36f_f0ef0665,
        64'h05130000_0517f87d,
        64'h959ff0ef_0ff00513,
        64'h347d4421_80826169,
        64'h6baa6b4a_6aea7a0a,
        64'h79aa794a_74ea640e,
        64'h852260ae_97dff0ef,
        64'h0ff00513_b09ff0ef,
        64'h45314581_46055479,
        64'hb7edf7ef_f0ef0ce5,
        64'h05130000_0517a809,
        64'h4401f520_4ee3197d,
        64'hc7910339_67b30347,
        64'h91638ade_93c117c2,
        64'h009567b3_9bdff0ef,
        64'h90c10ff0_051314c2,
        64'h0085149b_9cdff0ef,
        64'h0ff00513_fa9b93e3,
        64'h040a8a93_040b8b93,
        64'hfcda90e3_030a5a13,
        64'h06850307_9a138fb9,
        64'h00eb7733_0057171b,
        64'h0107571b_0107971b,
        64'h8fb900c7_971b8fb9,
        64'h8b3d0047_d71b8fb9,
        64'h93411742_01476733,
        64'h0006c783_008a5a1b,
        64'h008a171b_86dea9ff,
        64'hf0ef850a_04000593,
        64'h865e200b_8493040a,
        64'h8a934a01_8bd6fe85,
        64'h1ce3a43f_f0ef0ff0,
        64'h05133e80_09931b01,
        64'h0fe00413_6b090e05,
        64'h1b63bdff_f0ef4549,
        64'h4605fed7_9de307a1,
        64'h0114e398_577d878a,
        64'h02095913_8aaae55e,
        64'he95af152_f54efd26,
        64'he1a2e586_ed560206,
        64'h1913f94a_71558082,
        64'h91411542_8d3d8ff9,
        64'h17810057_171b6789,
        64'h0107571b_0105171b,
        64'h8d3d00c5_179b8d3d,
        64'h8bbd0045_579b00f5,
        64'hc53393c1_17c28fc9,
        64'h0085551b_0085179b,
        64'h808207f5_75138d3d,
        64'h0ff7f793_0045179b,
        64'h8d2d0ff5_75138d3d,
        64'h0045d51b_0075d79b,
        64'h8de9b7c5_5575b7d5,
        64'h55798082_6105557d,
        64'h690264a2_644260e2,
        64'h80826105_690264a2,
        64'h644260e2_4501c10d,
        64'heb9ff0ef_c115dd7f,
        64'hf0ef907f_f0efc4e5,
        64'h05130000_05179f3f,
        64'hf0ef4505_919ff0ef,
        64'h20850513_00000517,
        64'h925ff0ef_22450513,
        64'h00000517_931ff0ef,
        64'h21050513_00000517,
        64'hff2413e3_c8b9b57f,
        64'hf0ef0ff0_051334fd,
        64'h842ace7f_f0ef4501,
        64'h45810950_06134905,
        64'h71048493_6489f87d,
        64'hb79ff0ef_0ff00513,
        64'h347d4429_971ff0ef,
        64'h28850513_00000517,
        64'hafbff0ef_e04ae426,
        64'he822ec06_11018082,
        64'h61050015_351364a2,
        64'h64420004_051b60e2,
        64'hf69401e3_bb5ff0ef,
        64'h0ff00513_9a9ff0ef,
        64'hcf050513_00000517,
        64'ha95ff0ef_85229bbf,
        64'hf0ef2aa5_05130000,
        64'h05179c7f_f0ef2d65,
        64'h05130000_05179d3f,
        64'hf0ef2b25_05130000,
        64'h0517842a_d79ff0ef,
        64'h02900513_400005b7,
        64'h07700613_9f1ff0ef,
        64'hd3850513_00000517,
        64'haddff0ef_8522a03f,
        64'hf0ef2f25_05130000,
        64'h0517a0ff_f0ef3165,
        64'h05130000_0517a1bf,
        64'hf0ef2fa5_05130000,
        64'h0517c3bf_f0ef0ff0,
        64'h0513842a_dc9ff0ef,
        64'h03700513_45810650,
        64'h06134485_e822ec06,
        64'he4261101_80820141,
        64'h00153513_157d6402,
        64'h0004051b_60a2a5bf,
        64'hf0efda25_05130000,
        64'h0517b47f_f0ef8522,
        64'ha6dff0ef_35c50513,
        64'h00000517_a79ff0ef,
        64'h38050513_00000517,
        64'ha85ff0ef_36450513,
        64'h00000517_ca5ff0ef,
        64'h0ff00513_842ae33f,
        64'hf0efe022_e4060370,
        64'h05134581_06500613,
        64'h11418082_61050017,
        64'hb5136902_64a2f567,
        64'h87930009_079b6442,
        64'h60e2fe87_98e300f4,
        64'hf7938082_61056902,
        64'h64a26442_60e200f4,
        64'h08634501_4785cf7f,
        64'hf0ef0ff0_0513cfff,
        64'hf0ef0ff0_0513892a,
        64'hd09ff0ef_0ff00513,
        64'h84aad13f_f0ef0ff0,
        64'h0513d1bf_f0ef0ff0,
        64'h0513d23f_f0ef0ff0,
        64'h0513842a_eb1ff0ef,
        64'he04ae426_e822ec06,
        64'h45211aa0_05930870,
        64'h06131101_80826105,
        64'h45016902_64a26442,
        64'h60e28082_61054505,
        64'h690264a2_644260e2,
        64'hb4dff0ef_e9450513,
        64'h00000517_c39ff0ef,
        64'h4505b5ff_f0ef44e5,
        64'h05130000_0517b6bf,
        64'hf0ef46a5_05130000,
        64'h0517b77f_f0ef4565,
        64'h05130000_0517ff24,
        64'h13e3c4a9_d9dff0ef,
        64'h0ff00513_34fd842a,
        64'hf2dff0ef_45014581,
        64'h09500613_49057104,
        64'h8493e822_ec06e04a,
        64'h6489e426_1101be45,
        64'h6105efa5_05130000,
        64'h051764a2_60e26442,
        64'hca5ff0ef_8522bcbf,
        64'hf0ef4ba5_05130000,
        64'h0517bd7f_f0ef8526,
        64'hbddff0ef_842ee822,
        64'hec064c25_05130000,
        64'h051784aa_e4261101,
        64'h80826105_690264a2,
        64'h644260e2_fe07c6e3,
        64'h147d4187_d79b0185,
        64'h179be23f_f0ef0ff0,
        64'h0513cc01_a0110640,
        64'h0413e33f_f0ef8526,
        64'he39ff0ef_0ff47513,
        64'he41ff0ef_0ff57513,
        64'h0084551b_e4dff0ef,
        64'h0ff57513_0104551b,
        64'he59ff0ef_0184551b,
        64'he61ff0ef_04096513,
        64'he69ff0ef_84b2842e,
        64'he426e822_ec060ff0,
        64'h0513892a_e04a1101,
        64'hbdbd0ff0_05130030,
        64'h7032635f_30703264,
        64'h5f307032_665f3070,
        64'h32615f30_70326d5f,
        64'h30703269_34367672,
        64'h05100400_00002a01,
        64'h00766373_69720000,
        64'h00344100_203f3f79,
        64'h74706d65_20746f6e,
        64'h206f6669_66207872,
        64'h00000000_00000a0d,
        64'h2164657a_696c6169,
        64'h74696e69_20495053,
        64'h00000000_00007830,
        64'h203a7375_74617473,
        64'h00000000_00000a0d,
        64'h49505320_74696e69,
        64'h00008082_557dbf45,
        64'h47018082_4501d3b8,
        64'h4719dbb8_577d2000,
        64'h07b7fec7_19e3fef6,
        64'h0fa30605_55fcffe5,
        64'h8b8552fc_00c70b63,
        64'h200005b7_200006b7,
        64'h9732fff5_8b8552fc,
        64'h200006b7_d3b42000,
        64'h07b71060_0693fff5,
        64'h37fd0001_03200793,
        64'hfeb51ce3_d6bc0505,
        64'h00054783_200006b7,
        64'h00e505b3_93010205,
        64'h9713c5ad_dbb85779,
        64'h200007b7_06b7ed63,
        64'h10000793_b7d1d7bf,
        64'hf0ef0c25_05130000,
        64'h0517e19f_f0ef9101,
        64'h15025068_d91ff0ef,
        64'h0e050513_00000517,
        64'h80826105_64a20ff4,
        64'hf513d3b8_4719dbb8,
        64'h577d2000_07b76442,
        64'h60e2cf91_8b852481,
        64'h507c5464_fff58b85,
        64'h507c2000_0437d3b8,
        64'h10600713_200007b7,
        64'hfff537fd_00010640,
        64'h0793d7a8_dbb85779,
        64'he426e822_ec062000,
        64'h07b71101_b3fd6105,
        64'h12850513_00000517,
        64'h64a260e2_6442d03c,
        64'h4799e07f_f0ef14e5,
        64'h05130000_0517ea5f,
        64'hf0ef9101_02049513,
        64'h2481e1ff_f0ef1465,
        64'h05130000_05175064,
        64'hd03c1660_0793e33f,
        64'hf0ef17a5_05130000,
        64'h0517ed1f_f0ef9101,
        64'h02049513_2481e4bf,
        64'hf0ef1725_05130000,
        64'h05175064_d03c1040,
        64'h07932000_0437fff5,
        64'h37fd0001_47a9c3b8,
        64'h47292000_07b7e73f,
        64'hf0efe426_e822ec06,
        64'h19250513_11010000,
        64'h05178082_41088082,
        64'hc10c0000_30703263,
        64'h5f307032_645f3070,
        64'h32665f30_7032615f,
        64'h3070326d_5f307032,
        64'h69343676_72051004,
        64'h0000002a_01007663,
        64'h73697200_00003441,
        64'h00302e32_2e323120,
        64'h29672820_3a434347,
        64'h46454443_42413938,
        64'h37363534_33323130,
        64'h808200d7_0023dfe5,
        64'h0207f793_01474783,
        64'h10000737_00c70023,
        64'hdfe50207_f7930147,
        64'h47831000_07370007,
        64'h46830007_c60397aa,
        64'h973e8111_00f57713,
        64'h04078793_00000797,
        64'h8082fd16_15e33661,
        64'h01070023_dfe50207,
        64'hf7930147_478300d7,
        64'h0023dfe5_0207f793,
        64'h01474783_0006c683,
        64'h0007c803_96ae97ae,
        64'h8bbd8abd_0047d693,
        64'h00c557b3_58e11000,
        64'h073708e5_85930380,
        64'h06130000_05978082,
        64'hfd1615e3_36610107,
        64'h0023dfe5_0207f793,
        64'h01474783_00d70023,
        64'hdfe50207_f7930147,
        64'h47830006_c6830007,
        64'hc80396ae_97ae8bbd,
        64'h8abd0047_d69300c5,
        64'h57bb58e1_10000737,
        64'h0da58593_46610000,
        64'h05978082_00f58023,
        64'h0007c783_00e580a3,
        64'h97aa8111_00074703,
        64'h973e00f5_77130fe7,
        64'h87930000_07978082,
        64'hf6f50505_00154683,
        64'h00d70023_dfe50207,
        64'hf7930147_47831000,
        64'h0737ce91_00054683,
        64'h808200e7_88230200,
        64'h071300e7_8423fc70,
        64'h071300e7_8623470d,
        64'h00a78223_0ff57513,
        64'h00e78023_0085551b,
        64'h0ff57713_00e78623,
        64'hf8000713_00078223,
        64'h100007b7_02b5553b,
        64'h0045959b_808200a7,
        64'h0023dfe5_0207f793,
        64'h01474783_10000737,
        64'h80820205_75130147,
        64'hc5031000_07b78082,
        64'h00054503_808200b5,
        64'h0023000b_0a010800,
        64'h30703263_5f307032,
        64'h645f3070_32665f30,
        64'h7032615f_3070326d,
        64'h5f307032_69343676,
        64'h72050000_002c0100,
        64'h76637369_72000000,
        64'h36410032_2d746c75,
        64'h61666564_2d697274,
        64'h2c786e6c_7800746c,
        64'h75616665_642d6972,
        64'h742c786e_6c78006c,
        64'h6175642d_73692c78,
        64'h6e6c7800_746e6573,
        64'h6572702d_74707572,
        64'h7265746e_692c786e,
        64'h6c780068_74646977,
        64'h2d326f69_70672c78,
        64'h6e6c7800_68746469,
        64'h772d6f69_70672c78,
        64'h6e6c7800_322d746c,
        64'h75616665_642d7475,
        64'h6f642c78_6e6c7800,
        64'h746c7561_6665642d,
        64'h74756f64_2c786e6c,
        64'h7800322d_73747570,
        64'h6e692d6c_6c612c78,
        64'h6e6c7800_73747570,
        64'h6e692d6c_6c612c78,
        64'h6e6c7800_72656c6c,
        64'h6f72746e_6f632d6f,
        64'h69706700_736c6c65,
        64'h632d6f69_70672300,
        64'h73736572_6464612d,
        64'h63616d2d_6c61636f,
        64'h6c007077_2d656c62,
        64'h61736964_00736567,
        64'h6e61722d_65676174,
        64'h6c6f7600_79636e65,
        64'h75716572_662d7861,
        64'h6d2d6970_73006f69,
        64'h7461722d_6b63732c,
        64'h786e6c78_00737469,
        64'h622d7265_66736e61,
        64'h72742d6d_756e2c78,
        64'h6e6c7800_73746962,
        64'h2d73732d_6d756e2c,
        64'h786e6c78_00747369,
        64'h78652d6f_6669662c,
        64'h786e6c78_00796c69,
        64'h6d61662c_786e6c78,
        64'h00687464_69772d6f,
        64'h692d6765_72007466,
        64'h6968732d_67657200,
        64'h73747075_72726574,
        64'h6e690074_6e657261,
        64'h702d7470_75727265,
        64'h746e6900_64656570,
        64'h732d746e_65727275,
        64'h63007665_646e2c76,
        64'h63736972_00797469,
        64'h726f6972_702d7861,
        64'h6d2c7663_73697200,
        64'h73656d61_6e2d6765,
        64'h72006465_646e6574,
        64'h78652d73_74707572,
        64'h7265746e_69007365,
        64'h676e6172_00646564,
        64'h6e657073_75732d65,
        64'h74617473_2d6e6961,
        64'h74657200_72656767,
        64'h6972742d_746c7561,
        64'h6665642c_78756e69,
        64'h6c00736f_69706700,
        64'h656c646e_61687000,
        64'h72656c6c_6f72746e,
        64'h6f632d74_70757272,
        64'h65746e69_00736c6c,
        64'h65632d74_70757272,
        64'h65746e69_23007469,
        64'h6c70732d_626c7400,
        64'h65707974_2d756d6d,
        64'h00617369_2c766373,
        64'h69720073_75746174,
        64'h73006765_72006570,
        64'h79745f65_63697665,
        64'h64007963_6e657571,
        64'h6572662d_6b636f6c,
        64'h63007963_6e657571,
        64'h6572662d_65736162,
        64'h656d6974_00687461,
        64'h702d7475_6f647473,
        64'h006c6564_6f6d0065,
        64'h6c626974_61706d6f,
        64'h6300736c_6c65632d,
        64'h657a6973_2300736c,
        64'h6c65632d_73736572,
        64'h64646123_09000000,
        64'h02000000_02000000,
        64'h02000000_01000000,
        64'hb5000000_04000000,
        64'h03000000_ffffffff,
        64'hbf020000_04000000,
        64'h03000000_ffffffff,
        64'hae020000_04000000,
        64'h03000000_01000000,
        64'ha1020000_04000000,
        64'h03000000_00000000,
        64'h8a020000_04000000,
        64'h03000000_08000000,
        64'h79020000_04000000,
        64'h03000000_08000000,
        64'h69020000_04000000,
        64'h03000000_00000000,
        64'h55020000_04000000,
        64'h03000000_00000000,
        64'h43020000_04000000,
        64'h03000000_00000000,
        64'h31020000_04000000,
        64'h03000000_00000000,
        64'h21020000_04000000,
        64'h03000000_00000100,
        64'h00000000_00000040,
        64'h00000000_67000000,
        64'h10000000_03000000,
        64'h11020000_00000000,
        64'h03000000_00000000,
        64'h612e3030_2e312d6f,
        64'h6970672d_7370782c,
        64'h786e6c78_1b000000,
        64'h15000000_03000000,
        64'h02000000_05020000,
        64'h04000000_03000000,
        64'h00000030_30303030,
        64'h30303440_6f697067,
        64'h01000000_02000000,
        64'h00800000_00000000,
        64'h00000030_00000000,
        64'h67000000_10000000,
        64'h03000000_00007fe3,
        64'h023e1800_f3010000,
        64'h06000000_03000000,
        64'h00000000_03000000,
        64'h52010000_08000000,
        64'h03000000_03000000,
        64'h41010000_04000000,
        64'h03000000_006b726f,
        64'h7774656e_5b000000,
        64'h08000000_03000000,
        64'h00687465_2d637369,
        64'h72776f6c_1b000000,
        64'h0c000000_03000000,
        64'h00000000_30303030,
        64'h30303033_40687465,
        64'h2d637369_72776f6c,
        64'h01000000_02000000,
        64'h02000000_e8010000,
        64'h00000000_03000000,
        64'he40c0000_e40c0000,
        64'hd9010000_08000000,
        64'h03000000_20bcbe00,
        64'hc7010000_04000000,
        64'h03000000_00000000,
        64'h67000000_04000000,
        64'h03000000_00000000,
        64'h746f6c73_2d697073,
        64'h2d636d6d_1b000000,
        64'h0d000000_03000000,
        64'h00000030_40636d6d,
        64'h01000000_04000000,
        64'hb8010000_04000000,
        64'h03000000_08000000,
        64'ha1010000_04000000,
        64'h03000000_01000000,
        64'h90010000_04000000,
        64'h03000000_01000000,
        64'h80010000_04000000,
        64'h03000000_00003778,
        64'h69727461_74010000,
        64'h07000000_03000000,
        64'h00100000_00000000,
        64'h00000020_00000000,
        64'h67000000_10000000,
        64'h03000000_02000000,
        64'h02000000_52010000,
        64'h08000000_03000000,
        64'h03000000_41010000,
        64'h04000000_03000000,
        64'h00000000_0f000000,
        64'h04000000_03000000,
        64'h01000000_00000000,
        64'h04000000_03000000,
        64'h00612e30_302e322d,
        64'h6970732d_7370782c,
        64'h786e6c78_00622e30,
        64'h302e322d_6970732d,
        64'h7370782c_786e6c78,
        64'h1b000000_28000000,
        64'h03000000_00000000,
        64'h30303030_30303032,
        64'h40697073_01000000,
        64'h02000000_006c6f72,
        64'h746e6f63_0b010000,
        64'h08000000_03000000,
        64'h03000000_41010000,
        64'h04000000_03000000,
        64'h00100000_00000000,
        64'h00000018_00000000,
        64'h67000000_10000000,
        64'h03000000_07000000,
        64'h06000000_05000000,
        64'h04000000_52010000,
        64'h10000000_03000000,
        64'h00007265_6d69745f,
        64'h6270612c_706c7570,
        64'h1b000000_0f000000,
        64'h03000000_00003030,
        64'h30303030_38314072,
        64'h656d6974_01000000,
        64'h02000000_04000000,
        64'h67010000_04000000,
        64'h03000000_02000000,
        64'h5d010000_04000000,
        64'h03000000_01000000,
        64'h52010000_04000000,
        64'h03000000_03000000,
        64'h41010000_04000000,
        64'h03000000_00c20100,
        64'h33010000_04000000,
        64'h03000000_80f0fa02,
        64'h4b000000_04000000,
        64'h03000000_00100000,
        64'h00000000_00000010,
        64'h00000000_67000000,
        64'h10000000_03000000,
        64'h00000000_61303535,
        64'h3631736e_1b000000,
        64'h09000000_03000000,
        64'h00000030_30303030,
        64'h30303140_74726175,
        64'h01000000_02000000,
        64'h03000000_b5000000,
        64'h04000000_03000000,
        64'h1e000000_28010000,
        64'h04000000_03000000,
        64'h07000000_15010000,
        64'h04000000_03000000,
        64'h00000004_00000000,
        64'h0000000c_00000000,
        64'h67000000_10000000,
        64'h03000000_09000000,
        64'h02000000_0b000000,
        64'h02000000_f7000000,
        64'h10000000_03000000,
        64'ha0000000_00000000,
        64'h03000000_00306369,
        64'h6c702c76_63736972,
        64'h1b000000_0c000000,
        64'h03000000_01000000,
        64'h8f000000_04000000,
        64'h03000000_00000000,
        64'h00000000_04000000,
        64'h03000000_00000000,
        64'h30303030_30306340,
        64'h72656c6c_6f72746e,
        64'h6f632d74_70757272,
        64'h65746e69_01000000,
        64'h02000000_006c6f72,
        64'h746e6f63_0b010000,
        64'h08000000_03000000,
        64'h00000c00_00000000,
        64'h00000002_00000000,
        64'h67000000_10000000,
        64'h03000000_07000000,
        64'h02000000_03000000,
        64'h02000000_f7000000,
        64'h10000000_03000000,
        64'h00000000_30746e69,
        64'h6c632c76_63736972,
        64'h1b000000_0d000000,
        64'h03000000_00000030,
        64'h30303030_30324074,
        64'h6e696c63_01000000,
        64'hf0000000_00000000,
        64'h03000000_00007375,
        64'h622d656c_706d6973,
        64'h00636f73_2d657261,
        64'h622d656e_61697261,
        64'h2c687465_1b000000,
        64'h1f000000_03000000,
        64'h02000000_0f000000,
        64'h04000000_03000000,
        64'h02000000_00000000,
        64'h04000000_03000000,
        64'h00636f73_01000000,
        64'h02000000_02000000,
        64'hd9000000_00000000,
        64'h03000000_00000074,
        64'h61656274_72616568,
        64'hc3000000_0a000000,
        64'h03000000_00000000,
        64'h01000000_01000000,
        64'hbd000000_0c000000,
        64'h03000000_00000064,
        64'h656c2d74_61656274,
        64'h72616568_01000000,
        64'h00000073_64656c2d,
        64'h6f697067_1b000000,
        64'h0a000000_03000000,
        64'h00000000_7364656c,
        64'h01000000_02000000,
        64'h00000040_00000000,
        64'h00000080_00000000,
        64'h67000000_10000000,
        64'h03000000_00007972,
        64'h6f6d656d_5b000000,
        64'h07000000_03000000,
        64'h00303030_30303030,
        64'h38407972_6f6d656d,
        64'h01000000_02000000,
        64'h02000000_02000000,
        64'h02000000_b5000000,
        64'h04000000_03000000,
        64'h00006374_6e692d75,
        64'h70632c76_63736972,
        64'h1b000000_0f000000,
        64'h03000000_a0000000,
        64'h00000000_03000000,
        64'h01000000_8f000000,
        64'h04000000_03000000,
        64'h00000000_72656c6c,
        64'h6f72746e_6f632d74,
        64'h70757272_65746e69,
        64'h01000000_85000000,
        64'h00000000_03000000,
        64'h00003933_76732c76,
        64'h63736972_7c000000,
        64'h0b000000_03000000,
        64'h00000000_63616d69,
        64'h34367672_72000000,
        64'h09000000_03000000,
        64'h00000076_63736972,
        64'h00656e61_69726120,
        64'h2c687465_1b000000,
        64'h12000000_03000000,
        64'h00000000_79616b6f,
        64'h6b000000_05000000,
        64'h03000000_00000000,
        64'h67000000_04000000,
        64'h03000000_00757063,
        64'h5b000000_04000000,
        64'h03000000_80f0fa02,
        64'h4b000000_04000000,
        64'h03000000_00000030,
        64'h40757063_01000000,
        64'h40787d01_38000000,
        64'h04000000_03000000,
        64'h00000000_0f000000,
        64'h04000000_03000000,
        64'h01000000_00000000,
        64'h04000000_03000000,
        64'h00000000_73757063,
        64'h01000000_02000000,
        64'h00000030_30323531,
        64'h313a3030_30303030,
        64'h30314074_7261752f,
        64'h636f732f_2c000000,
        64'h1a000000_03000000,
        64'h00006e65_736f6863,
        64'h01000000_00657261,
        64'h622d656e_61697261,
        64'h2c687465_26000000,
        64'h10000000_03000000,
        64'h00766564_2d657261,
        64'h622d656e_61697261,
        64'h2c687465_1b000000,
        64'h14000000_03000000,
        64'h02000000_0f000000,
        64'h04000000_03000000,
        64'h02000000_00000000,
        64'h04000000_03000000,
        64'h00000000_01000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'he4080000_d2020000,
        64'h00000000_10000000,
        64'h11000000_28000000,
        64'h1c090000_38000000,
        64'hee0b0000_edfe0dd0,
        64'h00000000_00000000,
        64'h00008082_00000f93,
        64'h00000f13_00000e93,
        64'h00000e13_00000d93,
        64'h00000d13_00000c93,
        64'h00000c13_00000b93,
        64'h00000b13_00000a93,
        64'h00000a13_00000993,
        64'h00000913_00000893,
        64'h00000813_00000793,
        64'h00000713_00000693,
        64'h00000613_00000593,
        64'h00000513_00000493,
        64'h00000413_00000393,
        64'h00000313_00000293,
        64'h00000213_00000193,
        64'hb7cdfe03_0fe36322,
        64'h828202fe_0010029b,
        64'h09858593_00000597,
        64'hf1402573_020000ef,
        64'h0ff0000f_e4164285,
        64'hbfdd0321_00033023,
        64'h00230663_035a20f0,
        64'h031b5d50_e0ef0202,
        64'h9d63f140_22f3e402,
        64'h1141016a_0210011b
    };

    logic [$clog2(RomSize)-1:0] addr_q;

    always_ff @(posedge clk_i) begin
        if (req_i) begin
            addr_q <= addr_i[$clog2(RomSize)-1+3:3];
        end
    end

    // this prevents spurious Xes from propagating into
    // the speculative fetch stage of the core
    assign rdata_o = (addr_q < RomSize) ? mem[addr_q] : '0;
endmodule
